module data_inst(address, write_data, write, instruction, clk);

input clk;

input write;

input[31:0] write_data;

input[31:0] address;

output reg[0:31] instruction;//DATA INST sera a unica em EM BIG ENDIAN

//reg[0:31] registers[1000:0];//As instrucoes armazenadas tambem estao em BIG ENDIAN

wire[0:31] registers[1500:0];

/*always @(posedge clk)
begin	
	if(write)
	begin
		registers[address] <= write_data;
	end
end*/

always @(negedge clk)
begin
	instruction <= registers[address];
end


assign registers[0] = {32'b01110000000000000000000000000000};
assign registers[1] = {32'b10110001XXXXXXXXXXXXXXXXXXXXXXXX};
assign registers[2] = {32'b01111111000000000000000000000000};
assign registers[3] = {32'b01111101100000000000111111111111};
assign registers[4] = {32'b0110XXXX00000XXXXX11010000000001};
assign registers[5] = {32'b00010101110101101000000000000010};
assign registers[6] = {32'b1000000011010XXXXX11001XXXXXXXXX};
assign registers[7] = {32'b01000000000000000000000001110111};
assign registers[8] = {32'b0110XXXX11010XXXXX11001111111110};
assign registers[9] = {32'b0110XXXX11010XXXXX10100111111111};
assign registers[10] = {32'b0100001010100XXXXXXXXXXXXXXXXXXX};
assign registers[11] = {32'b00010101110111101100000000000001};
assign registers[12] = {32'b0110XXXX11011XXXXX01101000000000};
assign registers[13] = {32'b1010XXXX0110100000XXXX0000000000};
assign registers[14] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[15] = {32'b1000000000010XXXXX11000XXXXXXXXX};
assign registers[16] = {32'b00011000110000010111000XXXXXXXXX};
assign registers[17] = {32'b00010100110000001111000XXXXXXXXX};
assign registers[18] = {32'b00011000110000011111000XXXXXXXXX};
assign registers[19] = {32'b00010100110000010011000XXXXXXXXX};
assign registers[20] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[21] = {32'b1000000011111XXXXX01010XXXXXXXXX};
assign registers[22] = {32'b0110XXXX11011XXXXX00010000000011};
assign registers[23] = {32'b0110XXXX11011XXXXX00011000000010};
assign registers[24] = {32'b0110XXXX11011XXXXX00101000000001};
assign registers[25] = {32'b00010101110111101100000000000011};
assign registers[26] = {32'b01110010000000000000000000000001};
assign registers[27] = {32'b1000000000000XXXXX00110XXXXXXXXX};
assign registers[28] = {32'b1000000000101XXXXX00111XXXXXXXXX};
assign registers[29] = {32'b01110110100000000000000100000000};
assign registers[30] = {32'b01110111111111111111111111111111};
assign registers[31] = {32'b01000001000000000000000000001111};
assign registers[32] = {32'b1001XXXX0110011000XXXX0010000000};
assign registers[33] = {32'b01000011011000111100000000100111};
assign registers[34] = {32'b010100000011101100XXXXX000000001};
assign registers[35] = {32'b00010101001110011100000000000001};
assign registers[36] = {32'b00010101001100011000000000000001};
assign registers[37] = {32'b00010101110001100000000000000001};
assign registers[38] = {32'b01000000000000000000000000100000};
assign registers[39] = {32'b010100000010100110XXXXX000000000};
assign registers[40] = {32'b1000000000110XXXXX11000XXXXXXXXX};
assign registers[41] = {32'b0100001001010XXXXXXXXXXXXXXXXXXX};
assign registers[42] = {32'b0110XXXX11011XXXXX01100000000010};
assign registers[43] = {32'b0110XXXX11011XXXXX01101000000001};
assign registers[44] = {32'b00010101110111101100000000000010};
assign registers[45] = {32'b01110111000000000000000100000000};
assign registers[46] = {32'b0011XXXX0110001110XXXXXXXXXXXXXX};
assign registers[47] = {32'b10000001XXXXXXXXXX01111XXXXXXXXX};
assign registers[48] = {32'b010100000110101111XXXXX000000001};
assign registers[49] = {32'b10000010XXXXXXXXXX01100XXXXXXXXX};
assign registers[50] = {32'b0011XXXX0110001110XXXXXXXXXXXXXX};
assign registers[51] = {32'b10000001XXXXXXXXXX01111XXXXXXXXX};
assign registers[52] = {32'b010100000110101111XXXXX000000000};
assign registers[53] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[54] = {32'b0110XXXX11011XXXXX01100000001001};
assign registers[55] = {32'b0110XXXX11011XXXXX01101000001000};
assign registers[56] = {32'b01110111000000000000000000000111};
assign registers[57] = {32'b0010XXXX0110101110XXXXXXXXXXXXXX};
assign registers[58] = {32'b10000010XXXXXXXXXX01110XXXXXXXXX};
assign registers[59] = {32'b00010101011100111000000000000010};
assign registers[60] = {32'b00010100011100110001110XXXXXXXXX};
assign registers[61] = {32'b0110XXXX11011XXXXX01111000000111};
assign registers[62] = {32'b010100000111001111XXXXX000000000};
assign registers[63] = {32'b0110XXXX11011XXXXX01111000000110};
assign registers[64] = {32'b010100000111001111XXXXX000000001};
assign registers[65] = {32'b0110XXXX11011XXXXX01111000000101};
assign registers[66] = {32'b010100000111001111XXXXX000000010};
assign registers[67] = {32'b0110XXXX11011XXXXX01111000000100};
assign registers[68] = {32'b010100000111001111XXXXX000000011};
assign registers[69] = {32'b0110XXXX11011XXXXX01111000000011};
assign registers[70] = {32'b010100000111001111XXXXX000000100};
assign registers[71] = {32'b0110XXXX11011XXXXX01111000000010};
assign registers[72] = {32'b010100000111001111XXXXX000000101};
assign registers[73] = {32'b0110XXXX11011XXXXX01111000000001};
assign registers[74] = {32'b010100000111001111XXXXX000000110};
assign registers[75] = {32'b00010101110111101100000000001001};
assign registers[76] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[77] = {32'b0110XXXX11011XXXXX01100000000100};
assign registers[78] = {32'b0110XXXX11011XXXXX01101000000011};
assign registers[79] = {32'b0110XXXX11011XXXXX01110000000010};
assign registers[80] = {32'b0110XXXX11011XXXXX01111000000001};
assign registers[81] = {32'b00010101110111101100000000000100};
assign registers[82] = {32'b010100000110000000XXXXX000000000};
assign registers[83] = {32'b010100000110000000XXXXX000000001};
assign registers[84] = {32'b010100000110000000XXXXX000000010};
assign registers[85] = {32'b010100000110000000XXXXX000000011};
assign registers[86] = {32'b010100000110000000XXXXX000000100};
assign registers[87] = {32'b010100000110000000XXXXX000000101};
assign registers[88] = {32'b010100000110000000XXXXX000000110};
assign registers[89] = {32'b010100000110000000XXXXX000000111};
assign registers[90] = {32'b010100000110000000XXXXX000001000};
assign registers[91] = {32'b010100000110000000XXXXX000001001};
assign registers[92] = {32'b010100000110000000XXXXX000001010};
assign registers[93] = {32'b010100000110000000XXXXX000001011};
assign registers[94] = {32'b010100000110000000XXXXX000001100};
assign registers[95] = {32'b010100000110000000XXXXX000001101};
assign registers[96] = {32'b010100000110000000XXXXX000001110};
assign registers[97] = {32'b010100000110000000XXXXX000001111};
assign registers[98] = {32'b010100000110000000XXXXX000010000};
assign registers[99] = {32'b010100000110000000XXXXX000010001};
assign registers[100] = {32'b010100000110000000XXXXX000010010};
assign registers[101] = {32'b010100000110000000XXXXX000010011};
assign registers[102] = {32'b010100000110000000XXXXX000010100};
assign registers[103] = {32'b010100000110000000XXXXX000010101};
assign registers[104] = {32'b010100000110000000XXXXX000010110};
assign registers[105] = {32'b010100000110000000XXXXX000010111};
assign registers[106] = {32'b010100000110001101XXXXX000011000};
assign registers[107] = {32'b010100000110001110XXXXX000011001};
assign registers[108] = {32'b010100000110000000XXXXX000011010};
assign registers[109] = {32'b010100000110000000XXXXX000011011};
assign registers[110] = {32'b010100000110000000XXXXX000011100};
assign registers[111] = {32'b010100000110000000XXXXX000011101};
assign registers[112] = {32'b010100000110001111XXXXX000011110};
assign registers[113] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[114] = {32'b0110XXXX11011XXXXX11100000000011};
assign registers[115] = {32'b0110XXXX11011XXXXX11101000000010};
assign registers[116] = {32'b0110XXXX11011XXXXX00001000000001};
assign registers[117] = {32'b00010101110111101100000000000011};
assign registers[118] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[119] = {32'b1000000011001XXXXX11010XXXXXXXXX};
assign registers[120] = {32'b00010101110011100100000000010101};
assign registers[121] = {32'b00010101110011100100000001100100};
assign registers[122] = {32'b00010101110011100100000000000010};
assign registers[123] = {32'b01111010000000000000000001101110};
assign registers[124] = {32'b010100001101110100XXXXX000000000};
assign registers[125] = {32'b00010101110111101111111111111111};
assign registers[126] = {32'b010100001100100010XXXXX000000000};
assign registers[127] = {32'b010100001100100011XXXXX000000001};
assign registers[128] = {32'b010100001100100100XXXXX000000010};
assign registers[129] = {32'b010100001100100101XXXXX000000011};
assign registers[130] = {32'b010100001100100110XXXXX000000100};
assign registers[131] = {32'b010100001100100111XXXXX000000101};
assign registers[132] = {32'b010100001100101000XXXXX000000110};
assign registers[133] = {32'b010100001100101001XXXXX000000111};
assign registers[134] = {32'b010100001100101010XXXXX000001000};
assign registers[135] = {32'b00010101110011100100000000001001};
assign registers[136] = {32'b010100001100111010XXXXX000000000};
assign registers[137] = {32'b00010101110011100100000000000001};
assign registers[138] = {32'b01000001000000000000000000001011};
assign registers[139] = {32'b00010101110011100111111111111111};
assign registers[140] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[141] = {32'b00010101110011100111111111110111};
assign registers[142] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[143] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[144] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[145] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[146] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[147] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[148] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[149] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[150] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[151] = {32'b01111010000000000000000000000000};
assign registers[152] = {32'b01000011000101010000000010011010};
assign registers[153] = {32'b01000000000000000000001101101100};
assign registers[154] = {32'b01111010000000000000000000000001};
assign registers[155] = {32'b010100001101110100XXXXX000000000};
assign registers[156] = {32'b00010101110111101111111111111111};
assign registers[157] = {32'b01111010000000000000000000000000};
assign registers[158] = {32'b010100001101110100XXXXX000000000};
assign registers[159] = {32'b00010101110111101111111111111111};
assign registers[160] = {32'b01111010000000000000000000000000};
assign registers[161] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[162] = {32'b010100001101110100XXXXX000000000};
assign registers[163] = {32'b00010101110111101111111111111111};
assign registers[164] = {32'b010100001100100010XXXXX000000000};
assign registers[165] = {32'b010100001100100011XXXXX000000001};
assign registers[166] = {32'b010100001100100100XXXXX000000010};
assign registers[167] = {32'b010100001100100101XXXXX000000011};
assign registers[168] = {32'b010100001100100110XXXXX000000100};
assign registers[169] = {32'b010100001100100111XXXXX000000101};
assign registers[170] = {32'b010100001100101000XXXXX000000110};
assign registers[171] = {32'b010100001100101001XXXXX000000111};
assign registers[172] = {32'b010100001100101010XXXXX000001000};
assign registers[173] = {32'b00010101110011100100000000001001};
assign registers[174] = {32'b010100001100111010XXXXX000000000};
assign registers[175] = {32'b00010101110011100100000000000001};
assign registers[176] = {32'b01000001000000000000000000010101};
assign registers[177] = {32'b00010101110011100111111111111111};
assign registers[178] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[179] = {32'b00010101110011100111111111110111};
assign registers[180] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[181] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[182] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[183] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[184] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[185] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[186] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[187] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[188] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[189] = {32'b01111010000000000000000000000000};
assign registers[190] = {32'b01111010100000000000000000000000};
assign registers[191] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[192] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[193] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[194] = {32'b01111011000000000000000000000010};
assign registers[195] = {32'b00010100101011011001100XXXXXXXXX};
assign registers[196] = {32'b01111010000000000001000000000000};
assign registers[197] = {32'b0011XXXX1010001100XXXXXXXXXXXXXX};
assign registers[198] = {32'b10000010XXXXXXXXXX00100XXXXXXXXX};
assign registers[199] = {32'b01111010000000000000000000000000};
assign registers[200] = {32'b1000000010100XXXXX00011XXXXXXXXX};
assign registers[201] = {32'b1000000000100XXXXX00101XXXXXXXXX};
assign registers[202] = {32'b01111010000000000000000000000000};
assign registers[203] = {32'b01111010100000000000000000000000};
assign registers[204] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[205] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[206] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[207] = {32'b010100001101110101XXXXX000000000};
assign registers[208] = {32'b00010101110111101111111111111111};
assign registers[209] = {32'b010100001100100010XXXXX000000000};
assign registers[210] = {32'b010100001100100011XXXXX000000001};
assign registers[211] = {32'b010100001100100100XXXXX000000010};
assign registers[212] = {32'b010100001100100101XXXXX000000011};
assign registers[213] = {32'b010100001100100110XXXXX000000100};
assign registers[214] = {32'b010100001100100111XXXXX000000101};
assign registers[215] = {32'b010100001100101000XXXXX000000110};
assign registers[216] = {32'b010100001100101001XXXXX000000111};
assign registers[217] = {32'b010100001100101010XXXXX000001000};
assign registers[218] = {32'b00010101110011100100000000001001};
assign registers[219] = {32'b010100001100101100XXXXX000000000};
assign registers[220] = {32'b00010101110011100100000000000001};
assign registers[221] = {32'b010100001100111010XXXXX000000000};
assign registers[222] = {32'b00010101110011100100000000000001};
assign registers[223] = {32'b01000001000000000000000000001011};
assign registers[224] = {32'b00010101110011100111111111111111};
assign registers[225] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[226] = {32'b00010101110011100111111111111111};
assign registers[227] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[228] = {32'b00010101110011100111111111110111};
assign registers[229] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[230] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[231] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[232] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[233] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[234] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[235] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[236] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[237] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[238] = {32'b01111010000000000000000000000000};
assign registers[239] = {32'b01111010100000000000000000000000};
assign registers[240] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[241] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[242] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[243] = {32'b01000101000111010100000011110101};
assign registers[244] = {32'b01000000000000000000001101100011};
assign registers[245] = {32'b010100001101100011XXXXX000000000};
assign registers[246] = {32'b00010101110111101111111111111111};
assign registers[247] = {32'b010100001100100010XXXXX000000000};
assign registers[248] = {32'b010100001100100011XXXXX000000001};
assign registers[249] = {32'b010100001100100100XXXXX000000010};
assign registers[250] = {32'b010100001100100101XXXXX000000011};
assign registers[251] = {32'b010100001100100110XXXXX000000100};
assign registers[252] = {32'b010100001100100111XXXXX000000101};
assign registers[253] = {32'b010100001100101000XXXXX000000110};
assign registers[254] = {32'b010100001100101001XXXXX000000111};
assign registers[255] = {32'b010100001100101010XXXXX000001000};
assign registers[256] = {32'b00010101110011100100000000001001};
assign registers[257] = {32'b010100001100101100XXXXX000000000};
assign registers[258] = {32'b00010101110011100100000000000001};
assign registers[259] = {32'b010100001100111010XXXXX000000000};
assign registers[260] = {32'b00010101110011100100000000000001};
assign registers[261] = {32'b01000001000000000000000000001011};
assign registers[262] = {32'b00010101110011100111111111111111};
assign registers[263] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[264] = {32'b00010101110011100111111111111111};
assign registers[265] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[266] = {32'b00010101110011100111111111110111};
assign registers[267] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[268] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[269] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[270] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[271] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[272] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[273] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[274] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[275] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[276] = {32'b00010100001010010000110XXXXXXXXX};
assign registers[277] = {32'b01111010000000000000000000000001};
assign registers[278] = {32'b00010110001101010000110XXXXXXXXX};
assign registers[279] = {32'b01111010000000000000000000000001};
assign registers[280] = {32'b00010100000111010001101XXXXXXXXX};
assign registers[281] = {32'b01111010000000000000000000000000};
assign registers[282] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[283] = {32'b00010100101000110110100XXXXXXXXX};
assign registers[284] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[285] = {32'b010100001101110100XXXXX000000000};
assign registers[286] = {32'b00010101110111101111111111111111};
assign registers[287] = {32'b01111010000000000000000001111001};
assign registers[288] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[289] = {32'b010100001101110100XXXXX000000000};
assign registers[290] = {32'b00010101110111101111111111111111};
assign registers[291] = {32'b010100001100100010XXXXX000000000};
assign registers[292] = {32'b010100001100100011XXXXX000000001};
assign registers[293] = {32'b010100001100100100XXXXX000000010};
assign registers[294] = {32'b010100001100100101XXXXX000000011};
assign registers[295] = {32'b010100001100100110XXXXX000000100};
assign registers[296] = {32'b010100001100100111XXXXX000000101};
assign registers[297] = {32'b010100001100101000XXXXX000000110};
assign registers[298] = {32'b010100001100101001XXXXX000000111};
assign registers[299] = {32'b010100001100101010XXXXX000001000};
assign registers[300] = {32'b00010101110011100100000000001001};
assign registers[301] = {32'b010100001100101100XXXXX000000000};
assign registers[302] = {32'b010100001100101101XXXXX000000001};
assign registers[303] = {32'b00010101110011100100000000000010};
assign registers[304] = {32'b010100001100111010XXXXX000000000};
assign registers[305] = {32'b00010101110011100100000000000001};
assign registers[306] = {32'b01000001000000000000000000101010};
assign registers[307] = {32'b00010101110011100111111111111111};
assign registers[308] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[309] = {32'b00010101110011100111111111111110};
assign registers[310] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[311] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[312] = {32'b00010101110011100111111111110111};
assign registers[313] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[314] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[315] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[316] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[317] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[318] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[319] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[320] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[321] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[322] = {32'b01111010000000000000000000000000};
assign registers[323] = {32'b01111010100000000000000001111001};
assign registers[324] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[325] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[326] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[327] = {32'b010100001101110101XXXXX000000000};
assign registers[328] = {32'b00010101110111101111111111111111};
assign registers[329] = {32'b010100001100100010XXXXX000000000};
assign registers[330] = {32'b010100001100100011XXXXX000000001};
assign registers[331] = {32'b010100001100100100XXXXX000000010};
assign registers[332] = {32'b010100001100100101XXXXX000000011};
assign registers[333] = {32'b010100001100100110XXXXX000000100};
assign registers[334] = {32'b010100001100100111XXXXX000000101};
assign registers[335] = {32'b010100001100101000XXXXX000000110};
assign registers[336] = {32'b010100001100101001XXXXX000000111};
assign registers[337] = {32'b010100001100101010XXXXX000001000};
assign registers[338] = {32'b00010101110011100100000000001001};
assign registers[339] = {32'b010100001100101100XXXXX000000000};
assign registers[340] = {32'b010100001100101101XXXXX000000001};
assign registers[341] = {32'b00010101110011100100000000000010};
assign registers[342] = {32'b010100001100111010XXXXX000000000};
assign registers[343] = {32'b00010101110011100100000000000001};
assign registers[344] = {32'b01000001000000000000000000001011};
assign registers[345] = {32'b00010101110011100111111111111111};
assign registers[346] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[347] = {32'b00010101110011100111111111111110};
assign registers[348] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[349] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[350] = {32'b00010101110011100111111111110111};
assign registers[351] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[352] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[353] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[354] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[355] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[356] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[357] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[358] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[359] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[360] = {32'b01111010000000000000000000000001};
assign registers[361] = {32'b01111010100000000000000001111001};
assign registers[362] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[363] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[364] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[365] = {32'b010100001101110101XXXXX000000000};
assign registers[366] = {32'b00010101110111101111111111111111};
assign registers[367] = {32'b010100001100100010XXXXX000000000};
assign registers[368] = {32'b010100001100100011XXXXX000000001};
assign registers[369] = {32'b010100001100100100XXXXX000000010};
assign registers[370] = {32'b010100001100100101XXXXX000000011};
assign registers[371] = {32'b010100001100100110XXXXX000000100};
assign registers[372] = {32'b010100001100100111XXXXX000000101};
assign registers[373] = {32'b010100001100101000XXXXX000000110};
assign registers[374] = {32'b010100001100101001XXXXX000000111};
assign registers[375] = {32'b010100001100101010XXXXX000001000};
assign registers[376] = {32'b00010101110011100100000000001001};
assign registers[377] = {32'b010100001100101100XXXXX000000000};
assign registers[378] = {32'b010100001100101101XXXXX000000001};
assign registers[379] = {32'b00010101110011100100000000000010};
assign registers[380] = {32'b010100001100111010XXXXX000000000};
assign registers[381] = {32'b00010101110011100100000000000001};
assign registers[382] = {32'b01000001000000000000000000001011};
assign registers[383] = {32'b00010101110011100111111111111111};
assign registers[384] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[385] = {32'b00010101110011100111111111111110};
assign registers[386] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[387] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[388] = {32'b00010101110011100111111111110111};
assign registers[389] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[390] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[391] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[392] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[393] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[394] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[395] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[396] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[397] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[398] = {32'b01111010000000000000000000000000};
assign registers[399] = {32'b01111010100000000000000001111001};
assign registers[400] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[401] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[402] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[403] = {32'b010100001101110101XXXXX000000000};
assign registers[404] = {32'b00010101110111101111111111111111};
assign registers[405] = {32'b01111010000000000000000000000001};
assign registers[406] = {32'b01111010100000000000000001111001};
assign registers[407] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[408] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[409] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[410] = {32'b010100001101110101XXXXX000000000};
assign registers[411] = {32'b00010101110111101111111111111111};
assign registers[412] = {32'b010100001101100101XXXXX000000000};
assign registers[413] = {32'b00010101110111101111111111111111};
assign registers[414] = {32'b010100001100100010XXXXX000000000};
assign registers[415] = {32'b010100001100100011XXXXX000000001};
assign registers[416] = {32'b010100001100100100XXXXX000000010};
assign registers[417] = {32'b010100001100100101XXXXX000000011};
assign registers[418] = {32'b010100001100100110XXXXX000000100};
assign registers[419] = {32'b010100001100100111XXXXX000000101};
assign registers[420] = {32'b010100001100101000XXXXX000000110};
assign registers[421] = {32'b010100001100101001XXXXX000000111};
assign registers[422] = {32'b010100001100101010XXXXX000001000};
assign registers[423] = {32'b00010101110011100100000000001001};
assign registers[424] = {32'b010100001100101100XXXXX000000000};
assign registers[425] = {32'b010100001100101101XXXXX000000001};
assign registers[426] = {32'b00010101110011100100000000000010};
assign registers[427] = {32'b010100001100111010XXXXX000000000};
assign registers[428] = {32'b00010101110011100100000000000001};
assign registers[429] = {32'b01000001000000000000000000010101};
assign registers[430] = {32'b00010101110011100111111111111111};
assign registers[431] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[432] = {32'b00010101110011100111111111111110};
assign registers[433] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[434] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[435] = {32'b00010101110011100111111111110111};
assign registers[436] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[437] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[438] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[439] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[440] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[441] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[442] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[443] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[444] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[445] = {32'b1000000011000XXXXX00111XXXXXXXXX};
assign registers[446] = {32'b010100001101100101XXXXX000000000};
assign registers[447] = {32'b00010101110111101111111111111111};
assign registers[448] = {32'b010100001100100010XXXXX000000000};
assign registers[449] = {32'b010100001100100011XXXXX000000001};
assign registers[450] = {32'b010100001100100100XXXXX000000010};
assign registers[451] = {32'b010100001100100101XXXXX000000011};
assign registers[452] = {32'b010100001100100110XXXXX000000100};
assign registers[453] = {32'b010100001100100111XXXXX000000101};
assign registers[454] = {32'b010100001100101000XXXXX000000110};
assign registers[455] = {32'b010100001100101001XXXXX000000111};
assign registers[456] = {32'b010100001100101010XXXXX000001000};
assign registers[457] = {32'b00010101110011100100000000001001};
assign registers[458] = {32'b010100001100101100XXXXX000000000};
assign registers[459] = {32'b010100001100101101XXXXX000000001};
assign registers[460] = {32'b00010101110011100100000000000010};
assign registers[461] = {32'b010100001100111010XXXXX000000000};
assign registers[462] = {32'b00010101110011100100000000000001};
assign registers[463] = {32'b01000001000000000000000000001011};
assign registers[464] = {32'b00010101110011100111111111111111};
assign registers[465] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[466] = {32'b00010101110011100111111111111110};
assign registers[467] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[468] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[469] = {32'b00010101110011100111111111110111};
assign registers[470] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[471] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[472] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[473] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[474] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[475] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[476] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[477] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[478] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[479] = {32'b010100001101100111XXXXX000000000};
assign registers[480] = {32'b00010101110111101111111111111111};
assign registers[481] = {32'b010100001100100010XXXXX000000000};
assign registers[482] = {32'b010100001100100011XXXXX000000001};
assign registers[483] = {32'b010100001100100100XXXXX000000010};
assign registers[484] = {32'b010100001100100101XXXXX000000011};
assign registers[485] = {32'b010100001100100110XXXXX000000100};
assign registers[486] = {32'b010100001100100111XXXXX000000101};
assign registers[487] = {32'b010100001100101000XXXXX000000110};
assign registers[488] = {32'b010100001100101001XXXXX000000111};
assign registers[489] = {32'b010100001100101010XXXXX000001000};
assign registers[490] = {32'b00010101110011100100000000001001};
assign registers[491] = {32'b010100001100101100XXXXX000000000};
assign registers[492] = {32'b010100001100101101XXXXX000000001};
assign registers[493] = {32'b00010101110011100100000000000010};
assign registers[494] = {32'b010100001100111010XXXXX000000000};
assign registers[495] = {32'b00010101110011100100000000000001};
assign registers[496] = {32'b01000001000000000000000000001011};
assign registers[497] = {32'b00010101110011100111111111111111};
assign registers[498] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[499] = {32'b00010101110011100111111111111110};
assign registers[500] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[501] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[502] = {32'b00010101110011100111111111110111};
assign registers[503] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[504] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[505] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[506] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[507] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[508] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[509] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[510] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[511] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[512] = {32'b01111010000000000000000000000001};
assign registers[513] = {32'b00010100001011010001000XXXXXXXXX};
assign registers[514] = {32'b010100001101101000XXXXX000000000};
assign registers[515] = {32'b00010101110111101111111111111111};
assign registers[516] = {32'b010100001100100010XXXXX000000000};
assign registers[517] = {32'b010100001100100011XXXXX000000001};
assign registers[518] = {32'b010100001100100100XXXXX000000010};
assign registers[519] = {32'b010100001100100101XXXXX000000011};
assign registers[520] = {32'b010100001100100110XXXXX000000100};
assign registers[521] = {32'b010100001100100111XXXXX000000101};
assign registers[522] = {32'b010100001100101000XXXXX000000110};
assign registers[523] = {32'b010100001100101001XXXXX000000111};
assign registers[524] = {32'b010100001100101010XXXXX000001000};
assign registers[525] = {32'b00010101110011100100000000001001};
assign registers[526] = {32'b010100001100101100XXXXX000000000};
assign registers[527] = {32'b010100001100101101XXXXX000000001};
assign registers[528] = {32'b00010101110011100100000000000010};
assign registers[529] = {32'b010100001100111010XXXXX000000000};
assign registers[530] = {32'b00010101110011100100000000000001};
assign registers[531] = {32'b01000001000000000000000000001011};
assign registers[532] = {32'b00010101110011100111111111111111};
assign registers[533] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[534] = {32'b00010101110011100111111111111110};
assign registers[535] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[536] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[537] = {32'b00010101110011100111111111110111};
assign registers[538] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[539] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[540] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[541] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[542] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[543] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[544] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[545] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[546] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[547] = {32'b00010100010000011101001XXXXXXXXX};
assign registers[548] = {32'b01111010000000000000000000101000};
assign registers[549] = {32'b00010100010011010001010XXXXXXXXX};
assign registers[550] = {32'b010100001101100011XXXXX000000000};
assign registers[551] = {32'b00010101110111101111111111111111};
assign registers[552] = {32'b010100001100100010XXXXX000000000};
assign registers[553] = {32'b010100001100100011XXXXX000000001};
assign registers[554] = {32'b010100001100100100XXXXX000000010};
assign registers[555] = {32'b010100001100100101XXXXX000000011};
assign registers[556] = {32'b010100001100100110XXXXX000000100};
assign registers[557] = {32'b010100001100100111XXXXX000000101};
assign registers[558] = {32'b010100001100101000XXXXX000000110};
assign registers[559] = {32'b010100001100101001XXXXX000000111};
assign registers[560] = {32'b010100001100101010XXXXX000001000};
assign registers[561] = {32'b00010101110011100100000000001001};
assign registers[562] = {32'b010100001100101100XXXXX000000000};
assign registers[563] = {32'b010100001100101101XXXXX000000001};
assign registers[564] = {32'b00010101110011100100000000000010};
assign registers[565] = {32'b010100001100111010XXXXX000000000};
assign registers[566] = {32'b00010101110011100100000000000001};
assign registers[567] = {32'b01000001000000000000000000001011};
assign registers[568] = {32'b00010101110011100111111111111111};
assign registers[569] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[570] = {32'b00010101110011100111111111111110};
assign registers[571] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[572] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[573] = {32'b00010101110011100111111111110111};
assign registers[574] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[575] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[576] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[577] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[578] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[579] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[580] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[581] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[582] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[583] = {32'b010100001101101000XXXXX000000000};
assign registers[584] = {32'b00010101110111101111111111111111};
assign registers[585] = {32'b010100001100100010XXXXX000000000};
assign registers[586] = {32'b010100001100100011XXXXX000000001};
assign registers[587] = {32'b010100001100100100XXXXX000000010};
assign registers[588] = {32'b010100001100100101XXXXX000000011};
assign registers[589] = {32'b010100001100100110XXXXX000000100};
assign registers[590] = {32'b010100001100100111XXXXX000000101};
assign registers[591] = {32'b010100001100101000XXXXX000000110};
assign registers[592] = {32'b010100001100101001XXXXX000000111};
assign registers[593] = {32'b010100001100101010XXXXX000001000};
assign registers[594] = {32'b00010101110011100100000000001001};
assign registers[595] = {32'b010100001100101100XXXXX000000000};
assign registers[596] = {32'b010100001100101101XXXXX000000001};
assign registers[597] = {32'b00010101110011100100000000000010};
assign registers[598] = {32'b010100001100111010XXXXX000000000};
assign registers[599] = {32'b00010101110011100100000000000001};
assign registers[600] = {32'b01000001000000000000000000001011};
assign registers[601] = {32'b00010101110011100111111111111111};
assign registers[602] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[603] = {32'b00010101110011100111111111111110};
assign registers[604] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[605] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[606] = {32'b00010101110011100111111111110111};
assign registers[607] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[608] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[609] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[610] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[611] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[612] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[613] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[614] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[615] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[616] = {32'b010100001101100111XXXXX000000000};
assign registers[617] = {32'b00010101110111101111111111111111};
assign registers[618] = {32'b010100001100100010XXXXX000000000};
assign registers[619] = {32'b010100001100100011XXXXX000000001};
assign registers[620] = {32'b010100001100100100XXXXX000000010};
assign registers[621] = {32'b010100001100100101XXXXX000000011};
assign registers[622] = {32'b010100001100100110XXXXX000000100};
assign registers[623] = {32'b010100001100100111XXXXX000000101};
assign registers[624] = {32'b010100001100101000XXXXX000000110};
assign registers[625] = {32'b010100001100101001XXXXX000000111};
assign registers[626] = {32'b010100001100101010XXXXX000001000};
assign registers[627] = {32'b00010101110011100100000000001001};
assign registers[628] = {32'b010100001100101100XXXXX000000000};
assign registers[629] = {32'b010100001100101101XXXXX000000001};
assign registers[630] = {32'b00010101110011100100000000000010};
assign registers[631] = {32'b010100001100111010XXXXX000000000};
assign registers[632] = {32'b00010101110011100100000000000001};
assign registers[633] = {32'b01000001000000000000000000001011};
assign registers[634] = {32'b00010101110011100111111111111111};
assign registers[635] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[636] = {32'b00010101110011100111111111111110};
assign registers[637] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[638] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[639] = {32'b00010101110011100111111111110111};
assign registers[640] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[641] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[642] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[643] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[644] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[645] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[646] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[647] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[648] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[649] = {32'b010100001101101001XXXXX000000000};
assign registers[650] = {32'b00010101110111101111111111111111};
assign registers[651] = {32'b010100001100100010XXXXX000000000};
assign registers[652] = {32'b010100001100100011XXXXX000000001};
assign registers[653] = {32'b010100001100100100XXXXX000000010};
assign registers[654] = {32'b010100001100100101XXXXX000000011};
assign registers[655] = {32'b010100001100100110XXXXX000000100};
assign registers[656] = {32'b010100001100100111XXXXX000000101};
assign registers[657] = {32'b010100001100101000XXXXX000000110};
assign registers[658] = {32'b010100001100101001XXXXX000000111};
assign registers[659] = {32'b010100001100101010XXXXX000001000};
assign registers[660] = {32'b00010101110011100100000000001001};
assign registers[661] = {32'b010100001100101100XXXXX000000000};
assign registers[662] = {32'b010100001100101101XXXXX000000001};
assign registers[663] = {32'b00010101110011100100000000000010};
assign registers[664] = {32'b010100001100111010XXXXX000000000};
assign registers[665] = {32'b00010101110011100100000000000001};
assign registers[666] = {32'b01000001000000000000000000001011};
assign registers[667] = {32'b00010101110011100111111111111111};
assign registers[668] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[669] = {32'b00010101110011100111111111111110};
assign registers[670] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[671] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[672] = {32'b00010101110011100111111111110111};
assign registers[673] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[674] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[675] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[676] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[677] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[678] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[679] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[680] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[681] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[682] = {32'b010100001101101010XXXXX000000000};
assign registers[683] = {32'b00010101110111101111111111111111};
assign registers[684] = {32'b010100001100100010XXXXX000000000};
assign registers[685] = {32'b010100001100100011XXXXX000000001};
assign registers[686] = {32'b010100001100100100XXXXX000000010};
assign registers[687] = {32'b010100001100100101XXXXX000000011};
assign registers[688] = {32'b010100001100100110XXXXX000000100};
assign registers[689] = {32'b010100001100100111XXXXX000000101};
assign registers[690] = {32'b010100001100101000XXXXX000000110};
assign registers[691] = {32'b010100001100101001XXXXX000000111};
assign registers[692] = {32'b010100001100101010XXXXX000001000};
assign registers[693] = {32'b00010101110011100100000000001001};
assign registers[694] = {32'b010100001100101100XXXXX000000000};
assign registers[695] = {32'b010100001100101101XXXXX000000001};
assign registers[696] = {32'b00010101110011100100000000000010};
assign registers[697] = {32'b010100001100111010XXXXX000000000};
assign registers[698] = {32'b00010101110011100100000000000001};
assign registers[699] = {32'b01000001000000000000000000001011};
assign registers[700] = {32'b00010101110011100111111111111111};
assign registers[701] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[702] = {32'b00010101110011100111111111111110};
assign registers[703] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[704] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[705] = {32'b00010101110011100111111111110111};
assign registers[706] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[707] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[708] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[709] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[710] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[711] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[712] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[713] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[714] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[715] = {32'b010100001101100110XXXXX000000000};
assign registers[716] = {32'b00010101110111101111111111111111};
assign registers[717] = {32'b010100001100100010XXXXX000000000};
assign registers[718] = {32'b010100001100100011XXXXX000000001};
assign registers[719] = {32'b010100001100100100XXXXX000000010};
assign registers[720] = {32'b010100001100100101XXXXX000000011};
assign registers[721] = {32'b010100001100100110XXXXX000000100};
assign registers[722] = {32'b010100001100100111XXXXX000000101};
assign registers[723] = {32'b010100001100101000XXXXX000000110};
assign registers[724] = {32'b010100001100101001XXXXX000000111};
assign registers[725] = {32'b010100001100101010XXXXX000001000};
assign registers[726] = {32'b00010101110011100100000000001001};
assign registers[727] = {32'b010100001100101100XXXXX000000000};
assign registers[728] = {32'b010100001100101101XXXXX000000001};
assign registers[729] = {32'b00010101110011100100000000000010};
assign registers[730] = {32'b010100001100111010XXXXX000000000};
assign registers[731] = {32'b00010101110011100100000000000001};
assign registers[732] = {32'b01000001000000000000000000001011};
assign registers[733] = {32'b00010101110011100111111111111111};
assign registers[734] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[735] = {32'b00010101110011100111111111111110};
assign registers[736] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[737] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[738] = {32'b00010101110011100111111111110111};
assign registers[739] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[740] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[741] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[742] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[743] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[744] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[745] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[746] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[747] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[748] = {32'b01111010000000000000000000010101};
assign registers[749] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[750] = {32'b010100001101110100XXXXX000000000};
assign registers[751] = {32'b00010101110111101111111111111111};
assign registers[752] = {32'b010100001101100011XXXXX000000000};
assign registers[753] = {32'b00010101110111101111111111111111};
assign registers[754] = {32'b01111010000000000000000000000001};
assign registers[755] = {32'b00010100000111010001110XXXXXXXXX};
assign registers[756] = {32'b010100001101101110XXXXX000000000};
assign registers[757] = {32'b00010101110111101111111111111111};
assign registers[758] = {32'b01111010000000000000000000000000};
assign registers[759] = {32'b010100001101110100XXXXX000000000};
assign registers[760] = {32'b00010101110111101111111111111111};
assign registers[761] = {32'b010100001101101000XXXXX000000000};
assign registers[762] = {32'b00010101110111101111111111111111};
assign registers[763] = {32'b010100001101100111XXXXX000000000};
assign registers[764] = {32'b00010101110111101111111111111111};
assign registers[765] = {32'b010100001101101001XXXXX000000000};
assign registers[766] = {32'b00010101110111101111111111111111};
assign registers[767] = {32'b010100001101101010XXXXX000000000};
assign registers[768] = {32'b00010101110111101111111111111111};
assign registers[769] = {32'b010100001101100110XXXXX000000000};
assign registers[770] = {32'b00010101110111101111111111111111};
assign registers[771] = {32'b010100001100100010XXXXX000000000};
assign registers[772] = {32'b010100001100100011XXXXX000000001};
assign registers[773] = {32'b010100001100100100XXXXX000000010};
assign registers[774] = {32'b010100001100100101XXXXX000000011};
assign registers[775] = {32'b010100001100100110XXXXX000000100};
assign registers[776] = {32'b010100001100100111XXXXX000000101};
assign registers[777] = {32'b010100001100101000XXXXX000000110};
assign registers[778] = {32'b010100001100101001XXXXX000000111};
assign registers[779] = {32'b010100001100101010XXXXX000001000};
assign registers[780] = {32'b00010101110011100100000000001001};
assign registers[781] = {32'b010100001100101100XXXXX000000000};
assign registers[782] = {32'b010100001100101101XXXXX000000001};
assign registers[783] = {32'b010100001100101110XXXXX000000010};
assign registers[784] = {32'b00010101110011100100000000000011};
assign registers[785] = {32'b010100001100111010XXXXX000000000};
assign registers[786] = {32'b00010101110011100100000000000001};
assign registers[787] = {32'b01000001000000000000000000110110};
assign registers[788] = {32'b00010101110011100111111111111111};
assign registers[789] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[790] = {32'b00010101110011100111111111111101};
assign registers[791] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[792] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[793] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[794] = {32'b00010101110011100111111111110111};
assign registers[795] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[796] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[797] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[798] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[799] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[800] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[801] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[802] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[803] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[804] = {32'b010100001101101001XXXXX000000000};
assign registers[805] = {32'b00010101110111101111111111111111};
assign registers[806] = {32'b010100001101101010XXXXX000000000};
assign registers[807] = {32'b00010101110111101111111111111111};
assign registers[808] = {32'b010100001101100110XXXXX000000000};
assign registers[809] = {32'b00010101110111101111111111111111};
assign registers[810] = {32'b01111010000000000000000000000001};
assign registers[811] = {32'b00010100000111010001111XXXXXXXXX};
assign registers[812] = {32'b010100001101101111XXXXX000000000};
assign registers[813] = {32'b00010101110111101111111111111111};
assign registers[814] = {32'b010100001100100010XXXXX000000000};
assign registers[815] = {32'b010100001100100011XXXXX000000001};
assign registers[816] = {32'b010100001100100100XXXXX000000010};
assign registers[817] = {32'b010100001100100101XXXXX000000011};
assign registers[818] = {32'b010100001100100110XXXXX000000100};
assign registers[819] = {32'b010100001100100111XXXXX000000101};
assign registers[820] = {32'b010100001100101000XXXXX000000110};
assign registers[821] = {32'b010100001100101001XXXXX000000111};
assign registers[822] = {32'b010100001100101010XXXXX000001000};
assign registers[823] = {32'b00010101110011100100000000001001};
assign registers[824] = {32'b010100001100101100XXXXX000000000};
assign registers[825] = {32'b010100001100101101XXXXX000000001};
assign registers[826] = {32'b010100001100101110XXXXX000000010};
assign registers[827] = {32'b010100001100101111XXXXX000000011};
assign registers[828] = {32'b00010101110011100100000000000100};
assign registers[829] = {32'b010100001100111010XXXXX000000000};
assign registers[830] = {32'b00010101110011100100000000000001};
assign registers[831] = {32'b01000001000000000000000001001101};
assign registers[832] = {32'b00010101110011100111111111111111};
assign registers[833] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[834] = {32'b00010101110011100111111111111100};
assign registers[835] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[836] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[837] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[838] = {32'b0110XXXX11001XXXXX01111000000011};
assign registers[839] = {32'b00010101110011100111111111110111};
assign registers[840] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[841] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[842] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[843] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[844] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[845] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[846] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[847] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[848] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[849] = {32'b01111010000000000000000000000001};
assign registers[850] = {32'b00010100000111010000011XXXXXXXXX};
assign registers[851] = {32'b01111010000000000000000000000001};
assign registers[852] = {32'b00010100001101010000101XXXXXXXXX};
assign registers[853] = {32'b01111010000000000000000000000001};
assign registers[854] = {32'b01111010100000000000000000010101};
assign registers[855] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[856] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[857] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[858] = {32'b1000000010101XXXXX01000XXXXXXXXX};
assign registers[859] = {32'b01111010100000000000000000000001};
assign registers[860] = {32'b00010100010001010110100XXXXXXXXX};
assign registers[861] = {32'b01111011000000000000000000010101};
assign registers[862] = {32'b00010100101101101010110XXXXXXXXX};
assign registers[863] = {32'b01111011100000000000000000000001};
assign registers[864] = {32'b00010100101101011110111XXXXXXXXX};
assign registers[865] = {32'b010100001011110100XXXXX000000000};
assign registers[866] = {32'b01000000000000000000000011101110};
assign registers[867] = {32'b01111010000000000000000000000000};
assign registers[868] = {32'b1000000010100XXXXX01000XXXXXXXXX};
assign registers[869] = {32'b01111010100000000000000000000001};
assign registers[870] = {32'b00010110010001010110100XXXXXXXXX};
assign registers[871] = {32'b01111011000000000000000000010101};
assign registers[872] = {32'b00010100101101101010110XXXXXXXXX};
assign registers[873] = {32'b01111011100000000000000000000000};
assign registers[874] = {32'b00010100101101011110111XXXXXXXXX};
assign registers[875] = {32'b010100001011110100XXXXX000000000};
assign registers[876] = {32'b01111010000000000000000000000001};
assign registers[877] = {32'b01111010100000000000000000010101};
assign registers[878] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[879] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[880] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[881] = {32'b1000000010101XXXXX00010XXXXXXXXX};
assign registers[882] = {32'b01111010000000000000000010001100};
assign registers[883] = {32'b010100001101110100XXXXX000000000};
assign registers[884] = {32'b00010101110111101111111111111111};
assign registers[885] = {32'b010100001100100010XXXXX000000000};
assign registers[886] = {32'b010100001100100011XXXXX000000001};
assign registers[887] = {32'b010100001100100100XXXXX000000010};
assign registers[888] = {32'b010100001100100101XXXXX000000011};
assign registers[889] = {32'b010100001100100110XXXXX000000100};
assign registers[890] = {32'b010100001100100111XXXXX000000101};
assign registers[891] = {32'b010100001100101000XXXXX000000110};
assign registers[892] = {32'b010100001100101001XXXXX000000111};
assign registers[893] = {32'b010100001100101010XXXXX000001000};
assign registers[894] = {32'b00010101110011100100000000001001};
assign registers[895] = {32'b010100001100101100XXXXX000000000};
assign registers[896] = {32'b010100001100101101XXXXX000000001};
assign registers[897] = {32'b010100001100101110XXXXX000000010};
assign registers[898] = {32'b010100001100101111XXXXX000000011};
assign registers[899] = {32'b00010101110011100100000000000100};
assign registers[900] = {32'b010100001100111010XXXXX000000000};
assign registers[901] = {32'b00010101110011100100000000000001};
assign registers[902] = {32'b01000001000000000000000000001011};
assign registers[903] = {32'b00010101110011100111111111111111};
assign registers[904] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[905] = {32'b00010101110011100111111111111100};
assign registers[906] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[907] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[908] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[909] = {32'b0110XXXX11001XXXXX01111000000011};
assign registers[910] = {32'b00010101110011100111111111110111};
assign registers[911] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[912] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[913] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[914] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[915] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[916] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[917] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[918] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[919] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[920] = {32'b01111010000000000000000000000000};
assign registers[921] = {32'b01111010100000000000000000010101};
assign registers[922] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[923] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[924] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[925] = {32'b01111011000000000000000000000001};
assign registers[926] = {32'b00010100101011011000011XXXXXXXXX};
assign registers[927] = {32'b01111010000000000000000000000111};
assign registers[928] = {32'b0010XXXX0001110100XXXXXXXXXXXXXX};
assign registers[929] = {32'b10000010XXXXXXXXXX10000XXXXXXXXX};
assign registers[930] = {32'b01111010000000000000000000000011};
assign registers[931] = {32'b00010100101001000001000XXXXXXXXX};
assign registers[932] = {32'b01111010000000000000000000010101};
assign registers[933] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[934] = {32'b00010100101000100010100XXXXXXXXX};
assign registers[935] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[936] = {32'b01111010100000000000000000000000};
assign registers[937] = {32'b01000100101001010100001110101011};
assign registers[938] = {32'b01000000000000000000001111011110};
assign registers[939] = {32'b010100001101100011XXXXX000000000};
assign registers[940] = {32'b00010101110111101111111111111111};
assign registers[941] = {32'b010100001100100010XXXXX000000000};
assign registers[942] = {32'b010100001100100011XXXXX000000001};
assign registers[943] = {32'b010100001100100100XXXXX000000010};
assign registers[944] = {32'b010100001100100101XXXXX000000011};
assign registers[945] = {32'b010100001100100110XXXXX000000100};
assign registers[946] = {32'b010100001100100111XXXXX000000101};
assign registers[947] = {32'b010100001100101000XXXXX000000110};
assign registers[948] = {32'b010100001100101001XXXXX000000111};
assign registers[949] = {32'b010100001100101010XXXXX000001000};
assign registers[950] = {32'b00010101110011100100000000001001};
assign registers[951] = {32'b010100001100101100XXXXX000000000};
assign registers[952] = {32'b010100001100101101XXXXX000000001};
assign registers[953] = {32'b010100001100101110XXXXX000000010};
assign registers[954] = {32'b010100001100101111XXXXX000000011};
assign registers[955] = {32'b010100001100110000XXXXX000000100};
assign registers[956] = {32'b00010101110011100100000000000101};
assign registers[957] = {32'b010100001100111010XXXXX000000000};
assign registers[958] = {32'b00010101110011100100000000000001};
assign registers[959] = {32'b01000001000000000000000000001011};
assign registers[960] = {32'b00010101110011100111111111111111};
assign registers[961] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[962] = {32'b00010101110011100111111111111011};
assign registers[963] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[964] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[965] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[966] = {32'b0110XXXX11001XXXXX01111000000011};
assign registers[967] = {32'b0110XXXX11001XXXXX10000000000100};
assign registers[968] = {32'b00010101110011100111111111110111};
assign registers[969] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[970] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[971] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[972] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[973] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[974] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[975] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[976] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[977] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[978] = {32'b01111010000000000000000000000001};
assign registers[979] = {32'b00010100000111010000011XXXXXXXXX};
assign registers[980] = {32'b01001000000110001000001111010110};
assign registers[981] = {32'b01000000000000000000001111011000};
assign registers[982] = {32'b01111010000000000000000000000000};
assign registers[983] = {32'b1000000010100XXXXX00011XXXXXXXXX};
assign registers[984] = {32'b01111010000000000000000000000111};
assign registers[985] = {32'b0010XXXX0001110100XXXXXXXXXXXXXX};
assign registers[986] = {32'b10000010XXXXXXXXXX10001XXXXXXXXX};
assign registers[987] = {32'b01111010000000000000000000000011};
assign registers[988] = {32'b00010100101001000101000XXXXXXXXX};
assign registers[989] = {32'b01000000000000000000001110100100};
assign registers[990] = {32'b01111010000000000000000010010110};
assign registers[991] = {32'b010100001101110100XXXXX000000000};
assign registers[992] = {32'b00010101110111101111111111111111};
assign registers[993] = {32'b010100001100100010XXXXX000000000};
assign registers[994] = {32'b010100001100100011XXXXX000000001};
assign registers[995] = {32'b010100001100100100XXXXX000000010};
assign registers[996] = {32'b010100001100100101XXXXX000000011};
assign registers[997] = {32'b010100001100100110XXXXX000000100};
assign registers[998] = {32'b010100001100100111XXXXX000000101};
assign registers[999] = {32'b010100001100101000XXXXX000000110};
assign registers[1000] = {32'b010100001100101001XXXXX000000111};
assign registers[1001] = {32'b010100001100101010XXXXX000001000};
assign registers[1002] = {32'b00010101110011100100000000001001};
assign registers[1003] = {32'b010100001100101100XXXXX000000000};
assign registers[1004] = {32'b010100001100101101XXXXX000000001};
assign registers[1005] = {32'b010100001100101110XXXXX000000010};
assign registers[1006] = {32'b010100001100101111XXXXX000000011};
assign registers[1007] = {32'b010100001100110000XXXXX000000100};
assign registers[1008] = {32'b010100001100110001XXXXX000000101};
assign registers[1009] = {32'b00010101110011100100000000000110};
assign registers[1010] = {32'b010100001100111010XXXXX000000000};
assign registers[1011] = {32'b00010101110011100100000000000001};
assign registers[1012] = {32'b01000001000000000000000000001011};
assign registers[1013] = {32'b00010101110011100111111111111111};
assign registers[1014] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[1015] = {32'b00010101110011100111111111111010};
assign registers[1016] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[1017] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[1018] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[1019] = {32'b0110XXXX11001XXXXX01111000000011};
assign registers[1020] = {32'b0110XXXX11001XXXXX10000000000100};
assign registers[1021] = {32'b0110XXXX11001XXXXX10001000000101};
assign registers[1022] = {32'b00010101110011100111111111110111};
assign registers[1023] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[1024] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[1025] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[1026] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[1027] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[1028] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[1029] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[1030] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[1031] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[1032] = {32'b01111010000000000000000000000001};
assign registers[1033] = {32'b00010100010001010001000XXXXXXXXX};
assign registers[1034] = {32'b01111010000000000000000000000001};
assign registers[1035] = {32'b00010100010001010001001XXXXXXXXX};
assign registers[1036] = {32'b01111010000000000000000000000001};
assign registers[1037] = {32'b00010100010011010001010XXXXXXXXX};
assign registers[1038] = {32'b01111010000000000000000000010101};
assign registers[1039] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[1040] = {32'b00010100101000100010100XXXXXXXXX};
assign registers[1041] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[1042] = {32'b010100001101110100XXXXX000000000};
assign registers[1043] = {32'b00010101110111101111111111111111};
assign registers[1044] = {32'b010100001100100010XXXXX000000000};
assign registers[1045] = {32'b010100001100100011XXXXX000000001};
assign registers[1046] = {32'b010100001100100100XXXXX000000010};
assign registers[1047] = {32'b010100001100100101XXXXX000000011};
assign registers[1048] = {32'b010100001100100110XXXXX000000100};
assign registers[1049] = {32'b010100001100100111XXXXX000000101};
assign registers[1050] = {32'b010100001100101000XXXXX000000110};
assign registers[1051] = {32'b010100001100101001XXXXX000000111};
assign registers[1052] = {32'b010100001100101010XXXXX000001000};
assign registers[1053] = {32'b00010101110011100100000000001001};
assign registers[1054] = {32'b010100001100101100XXXXX000000000};
assign registers[1055] = {32'b010100001100101101XXXXX000000001};
assign registers[1056] = {32'b010100001100101110XXXXX000000010};
assign registers[1057] = {32'b010100001100101111XXXXX000000011};
assign registers[1058] = {32'b010100001100110000XXXXX000000100};
assign registers[1059] = {32'b010100001100110001XXXXX000000101};
assign registers[1060] = {32'b00010101110011100100000000000110};
assign registers[1061] = {32'b010100001100111010XXXXX000000000};
assign registers[1062] = {32'b00010101110011100100000000000001};
assign registers[1063] = {32'b01000001000000000000000000001011};
assign registers[1064] = {32'b00010101110011100111111111111111};
assign registers[1065] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[1066] = {32'b00010101110011100111111111111010};
assign registers[1067] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[1068] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[1069] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[1070] = {32'b0110XXXX11001XXXXX01111000000011};
assign registers[1071] = {32'b0110XXXX11001XXXXX10000000000100};
assign registers[1072] = {32'b0110XXXX11001XXXXX10001000000101};
assign registers[1073] = {32'b00010101110011100111111111110111};
assign registers[1074] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[1075] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[1076] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[1077] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[1078] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[1079] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[1080] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[1081] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[1082] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[1083] = {32'b01111010000000000000000000010101};
assign registers[1084] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[1085] = {32'b00010100101000100110100XXXXXXXXX};
assign registers[1086] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[1087] = {32'b010100001101110100XXXXX000000000};
assign registers[1088] = {32'b00010101110111101111111111111111};
assign registers[1089] = {32'b010100001100100010XXXXX000000000};
assign registers[1090] = {32'b010100001100100011XXXXX000000001};
assign registers[1091] = {32'b010100001100100100XXXXX000000010};
assign registers[1092] = {32'b010100001100100101XXXXX000000011};
assign registers[1093] = {32'b010100001100100110XXXXX000000100};
assign registers[1094] = {32'b010100001100100111XXXXX000000101};
assign registers[1095] = {32'b010100001100101000XXXXX000000110};
assign registers[1096] = {32'b010100001100101001XXXXX000000111};
assign registers[1097] = {32'b010100001100101010XXXXX000001000};
assign registers[1098] = {32'b00010101110011100100000000001001};
assign registers[1099] = {32'b010100001100101100XXXXX000000000};
assign registers[1100] = {32'b010100001100101101XXXXX000000001};
assign registers[1101] = {32'b010100001100101110XXXXX000000010};
assign registers[1102] = {32'b010100001100101111XXXXX000000011};
assign registers[1103] = {32'b010100001100110000XXXXX000000100};
assign registers[1104] = {32'b010100001100110001XXXXX000000101};
assign registers[1105] = {32'b00010101110011100100000000000110};
assign registers[1106] = {32'b010100001100111010XXXXX000000000};
assign registers[1107] = {32'b00010101110011100100000000000001};
assign registers[1108] = {32'b01000001000000000000000000001011};
assign registers[1109] = {32'b00010101110011100111111111111111};
assign registers[1110] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[1111] = {32'b00010101110011100111111111111010};
assign registers[1112] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[1113] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[1114] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[1115] = {32'b0110XXXX11001XXXXX01111000000011};
assign registers[1116] = {32'b0110XXXX11001XXXXX10000000000100};
assign registers[1117] = {32'b0110XXXX11001XXXXX10001000000101};
assign registers[1118] = {32'b00010101110011100111111111110111};
assign registers[1119] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[1120] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[1121] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[1122] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[1123] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[1124] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[1125] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[1126] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[1127] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[1128] = {32'b01111010000000000000000000010101};
assign registers[1129] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[1130] = {32'b00010100101000101010100XXXXXXXXX};
assign registers[1131] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[1132] = {32'b010100001101110100XXXXX000000000};
assign registers[1133] = {32'b00010101110111101111111111111111};
assign registers[1134] = {32'b010100001100100010XXXXX000000000};
assign registers[1135] = {32'b010100001100100011XXXXX000000001};
assign registers[1136] = {32'b010100001100100100XXXXX000000010};
assign registers[1137] = {32'b010100001100100101XXXXX000000011};
assign registers[1138] = {32'b010100001100100110XXXXX000000100};
assign registers[1139] = {32'b010100001100100111XXXXX000000101};
assign registers[1140] = {32'b010100001100101000XXXXX000000110};
assign registers[1141] = {32'b010100001100101001XXXXX000000111};
assign registers[1142] = {32'b010100001100101010XXXXX000001000};
assign registers[1143] = {32'b00010101110011100100000000001001};
assign registers[1144] = {32'b010100001100101100XXXXX000000000};
assign registers[1145] = {32'b010100001100101101XXXXX000000001};
assign registers[1146] = {32'b010100001100101110XXXXX000000010};
assign registers[1147] = {32'b010100001100101111XXXXX000000011};
assign registers[1148] = {32'b010100001100110000XXXXX000000100};
assign registers[1149] = {32'b010100001100110001XXXXX000000101};
assign registers[1150] = {32'b00010101110011100100000000000110};
assign registers[1151] = {32'b010100001100111010XXXXX000000000};
assign registers[1152] = {32'b00010101110011100100000000000001};
assign registers[1153] = {32'b01000001000000000000000000001011};
assign registers[1154] = {32'b00010101110011100111111111111111};
assign registers[1155] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[1156] = {32'b00010101110011100111111111111010};
assign registers[1157] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[1158] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[1159] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[1160] = {32'b0110XXXX11001XXXXX01111000000011};
assign registers[1161] = {32'b0110XXXX11001XXXXX10000000000100};
assign registers[1162] = {32'b0110XXXX11001XXXXX10001000000101};
assign registers[1163] = {32'b00010101110011100111111111110111};
assign registers[1164] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[1165] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[1166] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[1167] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[1168] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[1169] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[1170] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[1171] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[1172] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[1173] = {32'b01111010000000000000000000010101};
assign registers[1174] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[1175] = {32'b00010100101000100010100XXXXXXXXX};
assign registers[1176] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[1177] = {32'b010100001101110100XXXXX000000000};
assign registers[1178] = {32'b00010101110111101111111111111111};
assign registers[1179] = {32'b01111010000000000000000000010101};
assign registers[1180] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[1181] = {32'b00010100101000100110100XXXXXXXXX};
assign registers[1182] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[1183] = {32'b010100001101110100XXXXX000000000};
assign registers[1184] = {32'b00010101110111101111111111111111};
assign registers[1185] = {32'b01111010000000000000000000010101};
assign registers[1186] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[1187] = {32'b00010100101000101010100XXXXXXXXX};
assign registers[1188] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[1189] = {32'b010100001101110100XXXXX000000000};
assign registers[1190] = {32'b00010101110111101111111111111111};
assign registers[1191] = {32'b010100001100100010XXXXX000000000};
assign registers[1192] = {32'b010100001100100011XXXXX000000001};
assign registers[1193] = {32'b010100001100100100XXXXX000000010};
assign registers[1194] = {32'b010100001100100101XXXXX000000011};
assign registers[1195] = {32'b010100001100100110XXXXX000000100};
assign registers[1196] = {32'b010100001100100111XXXXX000000101};
assign registers[1197] = {32'b010100001100101000XXXXX000000110};
assign registers[1198] = {32'b010100001100101001XXXXX000000111};
assign registers[1199] = {32'b010100001100101010XXXXX000001000};
assign registers[1200] = {32'b00010101110011100100000000001001};
assign registers[1201] = {32'b010100001100101100XXXXX000000000};
assign registers[1202] = {32'b010100001100101101XXXXX000000001};
assign registers[1203] = {32'b010100001100101110XXXXX000000010};
assign registers[1204] = {32'b010100001100101111XXXXX000000011};
assign registers[1205] = {32'b010100001100110000XXXXX000000100};
assign registers[1206] = {32'b010100001100110001XXXXX000000101};
assign registers[1207] = {32'b00010101110011100100000000000110};
assign registers[1208] = {32'b010100001100111010XXXXX000000000};
assign registers[1209] = {32'b00010101110011100100000000000001};
assign registers[1210] = {32'b01000001000000000000000001110010};
assign registers[1211] = {32'b00010101110011100111111111111111};
assign registers[1212] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[1213] = {32'b00010101110011100111111111111010};
assign registers[1214] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[1215] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[1216] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[1217] = {32'b0110XXXX11001XXXXX01111000000011};
assign registers[1218] = {32'b0110XXXX11001XXXXX10000000000100};
assign registers[1219] = {32'b0110XXXX11001XXXXX10001000000101};
assign registers[1220] = {32'b00010101110011100111111111110111};
assign registers[1221] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[1222] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[1223] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[1224] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[1225] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[1226] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[1227] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[1228] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[1229] = {32'b0110XXXX11001XXXXX01010000001000};
assign registers[1230] = {32'b10110010XXXXXXXXXXXXXXXXXXXXXXXX};
assign registers[1231] = {32'b00000001000000000000000000000000};
assign registers[1232] = {32'b11111111111111111111111111111111};

endmodule 