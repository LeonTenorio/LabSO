module disk_controller(
input[2:0] track,
input[4:0] sector,
input[6:0] address_in_sector,
input read,
input write,
input[31:0] write_value,
output reg[31:0] read_value,
output reg read_done,
output reg write_done,
input clk
);

reg[31:0] values[32768:0];
wire[31:0] registers[32768:0];
reg not_initial[32768:0];

reg not_first_clk = 0;

always @(posedge clk)
begin
	write_done = 0;
	if(write)
	begin
		values[{track, sector, address_in_sector}] = write_value;
		not_initial[{track, sector, address_in_sector}] = 1;
		write_done = 1;
	end
end

always @(negedge clk)
begin
	read_done = 0;
	if(read)
	begin
		if(not_initial[{track, sector, address_in_sector}])
		begin
			read_value = values[{track, sector, address_in_sector}];
		end
		else
		begin
			read_value = registers[{track, sector, address_in_sector}];
		end
		read_done = 1;
	end
end

assign registers[0] = {16'd0, 16'd696};
assign registers[1] = {32'd300};
assign registers[2] = {32'b01110000000000000000000000000000};
assign registers[3] = {32'b10110001XXXXXXXXXXXXXXXXXXXXXXXX};
assign registers[4] = {32'b01111111000000000000000000000000};
assign registers[5] = {32'b01111101100000000000111111111111};
assign registers[6] = {32'b0110XXXX00000XXXXX11010000000001};
assign registers[7] = {32'b00010101110101101000000000001010};
assign registers[8] = {32'b1000000011010XXXXX11001XXXXXXXXX};
assign registers[9] = {32'b01000000000000000000000001101001};
assign registers[10] = {32'b0110XXXX11010XXXXX11001111111110};
assign registers[11] = {32'b0110XXXX11010XXXXX10100111111111};
assign registers[12] = {32'b0100001010100XXXXXXXXXXXXXXXXXXX};
assign registers[13] = {32'b0110XXXX11011XXXXX00010000000010};
assign registers[14] = {32'b0110XXXX11011XXXXX00011000000001};
assign registers[15] = {32'b00010101110111101100000000000010};
assign registers[16] = {32'b00010101000110110000000000011011};
assign registers[17] = {32'b0110XXXX01100XXXXX01100000000000};
assign registers[18] = {32'b00010100011000001001100XXXXXXXXX};
assign registers[19] = {32'b0110XXXX01100XXXXX11000000000000};
assign registers[20] = {32'b00011001110001100011000XXXXXXXXX};
assign registers[21] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[22] = {32'b00010101110111101100000000000001};
assign registers[23] = {32'b0110XXXX11011XXXXX01101000000000};
assign registers[24] = {32'b1010XXXX0110100000XXXX0000000000};
assign registers[25] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[26] = {32'b1000000000010XXXXX11000XXXXXXXXX};
assign registers[27] = {32'b00011000110000010111000XXXXXXXXX};
assign registers[28] = {32'b00010100110000001111000XXXXXXXXX};
assign registers[29] = {32'b00011000110000011111000XXXXXXXXX};
assign registers[30] = {32'b00010100110000010011000XXXXXXXXX};
assign registers[31] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[32] = {32'b1000000011111XXXXX01010XXXXXXXXX};
assign registers[33] = {32'b0110XXXX11011XXXXX00010000000011};
assign registers[34] = {32'b0110XXXX11011XXXXX00011000000010};
assign registers[35] = {32'b0110XXXX11011XXXXX00101000000001};
assign registers[36] = {32'b00010101110111101100000000000011};
assign registers[37] = {32'b01110010000000000000000000000001};
assign registers[38] = {32'b1000000000000XXXXX00110XXXXXXXXX};
assign registers[39] = {32'b1000000000101XXXXX00111XXXXXXXXX};
assign registers[40] = {32'b01110110100000000000000100000000};
assign registers[41] = {32'b01110111111111111111111111111111};
assign registers[42] = {32'b01000001000000000000000000011000};
assign registers[43] = {32'b1001XXXX0110011000XXXX0010000000};
assign registers[44] = {32'b01000011011000111100000000110000};
assign registers[45] = {32'b010100000011101100XXXXX000000001};
assign registers[46] = {32'b00010101001110011100000000000001};
assign registers[47] = {32'b00010101001100011000000000000001};
assign registers[48] = {32'b00010101110001100000000000000001};
assign registers[49] = {32'b01000000000000000000000000101001};
assign registers[50] = {32'b010100000010100110XXXXX000000000};
assign registers[51] = {32'b1000000000110XXXXX11000XXXXXXXXX};
assign registers[52] = {32'b0100001001010XXXXXXXXXXXXXXXXXXX};
assign registers[53] = {32'b0110XXXX11011XXXXX01100000000010};
assign registers[54] = {32'b0110XXXX11011XXXXX01101000000001};
assign registers[55] = {32'b00010101110111101100000000000010};
assign registers[56] = {32'b01110111000000000000000100000000};
assign registers[57] = {32'b0011XXXX0110001110XXXXXXXXXXXXXX};
assign registers[58] = {32'b10000001XXXXXXXXXX01111XXXXXXXXX};
assign registers[59] = {32'b010100000110101111XXXXX000000001};
assign registers[60] = {32'b10000010XXXXXXXXXX01100XXXXXXXXX};
assign registers[61] = {32'b0011XXXX0110001110XXXXXXXXXXXXXX};
assign registers[62] = {32'b10000001XXXXXXXXXX01111XXXXXXXXX};
assign registers[63] = {32'b010100000110101111XXXXX000000000};
assign registers[64] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[65] = {32'b0110XXXX11011XXXXX01100000000100};
assign registers[66] = {32'b0110XXXX11011XXXXX01101000000011};
assign registers[67] = {32'b0110XXXX11011XXXXX01110000000010};
assign registers[68] = {32'b0110XXXX11011XXXXX01111000000001};
assign registers[69] = {32'b00010101110111101100000000000100};
assign registers[70] = {32'b010100000110000000XXXXX000000000};
assign registers[71] = {32'b010100000110000000XXXXX000000001};
assign registers[72] = {32'b010100000110000000XXXXX000000010};
assign registers[73] = {32'b010100000110000000XXXXX000000011};
assign registers[74] = {32'b010100000110000000XXXXX000000100};
assign registers[75] = {32'b010100000110000000XXXXX000000101};
assign registers[76] = {32'b010100000110000000XXXXX000000110};
assign registers[77] = {32'b010100000110000000XXXXX000000111};
assign registers[78] = {32'b010100000110000000XXXXX000001000};
assign registers[79] = {32'b010100000110000000XXXXX000001001};
assign registers[80] = {32'b010100000110000000XXXXX000001010};
assign registers[81] = {32'b010100000110000000XXXXX000001011};
assign registers[82] = {32'b010100000110000000XXXXX000001100};
assign registers[83] = {32'b010100000110000000XXXXX000001101};
assign registers[84] = {32'b010100000110000000XXXXX000001110};
assign registers[85] = {32'b010100000110000000XXXXX000001111};
assign registers[86] = {32'b010100000110000000XXXXX000010000};
assign registers[87] = {32'b010100000110000000XXXXX000010001};
assign registers[88] = {32'b010100000110000000XXXXX000010010};
assign registers[89] = {32'b010100000110000000XXXXX000010011};
assign registers[90] = {32'b010100000110000000XXXXX000010100};
assign registers[91] = {32'b010100000110000000XXXXX000010101};
assign registers[92] = {32'b010100000110000000XXXXX000010110};
assign registers[93] = {32'b010100000110001101XXXXX000010111};
assign registers[94] = {32'b010100000110001101XXXXX000011000};
assign registers[95] = {32'b010100000110001110XXXXX000011001};
assign registers[96] = {32'b010100000110000000XXXXX000011010};
assign registers[97] = {32'b010100000110000000XXXXX000011011};
assign registers[98] = {32'b010100000110000000XXXXX000011100};
assign registers[99] = {32'b010100000110000000XXXXX000011101};
assign registers[100] = {32'b010100000110001111XXXXX000011110};
assign registers[101] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[102] = {32'b0110XXXX11011XXXXX11100000000011};
assign registers[103] = {32'b0110XXXX11011XXXXX11101000000010};
assign registers[104] = {32'b0110XXXX11011XXXXX00001000000001};
assign registers[105] = {32'b00010101110111101100000000000011};
assign registers[106] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[107] = {32'b1000000011001XXXXX11010XXXXXXXXX};
assign registers[108] = {32'b00010101110011100100000000010101};
assign registers[109] = {32'b00010101110011100100000010001000};
assign registers[110] = {32'b00010101110011100100000000000010};
assign registers[111] = {32'b01111010000000000000000000000001};
assign registers[112] = {32'b01111010100000000000000000010101};
assign registers[113] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[114] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[115] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[116] = {32'b01111011000000000000000000000000};
assign registers[117] = {32'b01000100101011011000000001110101};
assign registers[118] = {32'b01000000000000000000000011011001};
assign registers[119] = {32'b01111010000000000000000000000000};
assign registers[120] = {32'b01111010100000000000000000010101};
assign registers[121] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[122] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[123] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[124] = {32'b1000000010101XXXXX00010XXXXXXXXX};
assign registers[125] = {32'b01111010000000000000000000000111};
assign registers[126] = {32'b0010XXXX1010000010XXXXXXXXXXXXXX};
assign registers[127] = {32'b10000010XXXXXXXXXX00111XXXXXXXXX};
assign registers[128] = {32'b01111010000000000000000000000101};
assign registers[129] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[130] = {32'b01111010000000000000000000000010};
assign registers[131] = {32'b00010100001111010001000XXXXXXXXX};
assign registers[132] = {32'b01111010000000000000000000010101};
assign registers[133] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[134] = {32'b00010100101000011110100XXXXXXXXX};
assign registers[135] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[136] = {32'b010100001101110100XXXXX000000000};
assign registers[137] = {32'b00010101110111101111111111111111};
assign registers[138] = {32'b01111010000000000000000000010101};
assign registers[139] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[140] = {32'b00010100101000100010100XXXXXXXXX};
assign registers[141] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[142] = {32'b010100001101110100XXXXX000000000};
assign registers[143] = {32'b00010101110111101111111111111111};
assign registers[144] = {32'b010100001100100010XXXXX000000000};
assign registers[145] = {32'b010100001100100011XXXXX000000001};
assign registers[146] = {32'b010100001100100100XXXXX000000010};
assign registers[147] = {32'b010100001100100101XXXXX000000011};
assign registers[148] = {32'b010100001100100110XXXXX000000100};
assign registers[149] = {32'b010100001100100111XXXXX000000101};
assign registers[150] = {32'b010100001100101000XXXXX000000110};
assign registers[151] = {32'b010100001100101001XXXXX000000111};
assign registers[152] = {32'b00010101110011100100000000001000};
assign registers[153] = {32'b010100001100111010XXXXX000000000};
assign registers[154] = {32'b00010101110011100100000000000001};
assign registers[155] = {32'b01000001000000000000000000001011};
assign registers[156] = {32'b00010101110011100111111111111111};
assign registers[157] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[158] = {32'b00010101110011100111111111111000};
assign registers[159] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[160] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[161] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[162] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[163] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[164] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[165] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[166] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[167] = {32'b1000000011000XXXXX01001XXXXXXXXX};
assign registers[168] = {32'b01111010000000000000000000000001};
assign registers[169] = {32'b01000011010011010000000010101001};
assign registers[170] = {32'b01000000000000000000000011011001};
assign registers[171] = {32'b01111010000000000000000010010110};
assign registers[172] = {32'b010100001101110100XXXXX000000000};
assign registers[173] = {32'b00010101110111101111111111111111};
assign registers[174] = {32'b010100001100100010XXXXX000000000};
assign registers[175] = {32'b010100001100100011XXXXX000000001};
assign registers[176] = {32'b010100001100100100XXXXX000000010};
assign registers[177] = {32'b010100001100100101XXXXX000000011};
assign registers[178] = {32'b010100001100100110XXXXX000000100};
assign registers[179] = {32'b010100001100100111XXXXX000000101};
assign registers[180] = {32'b010100001100101000XXXXX000000110};
assign registers[181] = {32'b010100001100101001XXXXX000000111};
assign registers[182] = {32'b00010101110011100100000000001000};
assign registers[183] = {32'b010100001100111010XXXXX000000000};
assign registers[184] = {32'b00010101110011100100000000000001};
assign registers[185] = {32'b01000001000000000000000000010100};
assign registers[186] = {32'b00010101110011100111111111111111};
assign registers[187] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[188] = {32'b00010101110011100111111111111000};
assign registers[189] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[190] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[191] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[192] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[193] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[194] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[195] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[196] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[197] = {32'b01111010000000000000000000000001};
assign registers[198] = {32'b00010110001111010000111XXXXXXXXX};
assign registers[199] = {32'b01111010000000000000000000000010};
assign registers[200] = {32'b1000000010100XXXXX10101XXXXXXXXX};
assign registers[201] = {32'b01111011000000000000000000010101};
assign registers[202] = {32'b00010100101101101010110XXXXXXXXX};
assign registers[203] = {32'b00010100101100011110111XXXXXXXXX};
assign registers[204] = {32'b010100001011110101XXXXX000000000};
assign registers[205] = {32'b01111010000000000000000000000001};
assign registers[206] = {32'b01111010100000000000000000010101};
assign registers[207] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[208] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[209] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[210] = {32'b1000000010101XXXXX00111XXXXXXXXX};
assign registers[211] = {32'b01111010000000000000000000000001};
assign registers[212] = {32'b00010110001111010000111XXXXXXXXX};
assign registers[213] = {32'b1000000000111XXXXX10100XXXXXXXXX};
assign registers[214] = {32'b01111010100000000000000000010101};
assign registers[215] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[216] = {32'b01111011000000000000000000000001};
assign registers[217] = {32'b00010100101011011010110XXXXXXXXX};
assign registers[218] = {32'b010100001011010100XXXXX000000000};
assign registers[219] = {32'b01111010000000000000000000000001};
assign registers[220] = {32'b01111010100000000000000000010101};
assign registers[221] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[222] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[223] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[224] = {32'b01111011000000000000000000000000};
assign registers[225] = {32'b01000011101011011000000011100001};
assign registers[226] = {32'b01000000000000000000001000100101};
assign registers[227] = {32'b01111010000000000000000000000001};
assign registers[228] = {32'b010100001101110100XXXXX000000000};
assign registers[229] = {32'b00010101110111101111111111111111};
assign registers[230] = {32'b01111010000000000000000000000000};
assign registers[231] = {32'b010100001101110100XXXXX000000000};
assign registers[232] = {32'b00010101110111101111111111111111};
assign registers[233] = {32'b01111010000000000000000000000000};
assign registers[234] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[235] = {32'b010100001101110100XXXXX000000000};
assign registers[236] = {32'b00010101110111101111111111111111};
assign registers[237] = {32'b010100001100100010XXXXX000000000};
assign registers[238] = {32'b010100001100100011XXXXX000000001};
assign registers[239] = {32'b010100001100100100XXXXX000000010};
assign registers[240] = {32'b010100001100100101XXXXX000000011};
assign registers[241] = {32'b010100001100100110XXXXX000000100};
assign registers[242] = {32'b010100001100100111XXXXX000000101};
assign registers[243] = {32'b010100001100101000XXXXX000000110};
assign registers[244] = {32'b010100001100101001XXXXX000000111};
assign registers[245] = {32'b00010101110011100100000000001000};
assign registers[246] = {32'b010100001100111010XXXXX000000000};
assign registers[247] = {32'b00010101110011100100000000000001};
assign registers[248] = {32'b01000001000000000000000000011110};
assign registers[249] = {32'b00010101110011100111111111111111};
assign registers[250] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[251] = {32'b00010101110011100111111111111000};
assign registers[252] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[253] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[254] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[255] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[256] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[257] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[258] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[259] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[260] = {32'b01111010000000000001000000000000};
assign registers[261] = {32'b1000000010100XXXXX00100XXXXXXXXX};
assign registers[262] = {32'b01111010000000000000000010011101};
assign registers[263] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[264] = {32'b00010110001001010000100XXXXXXXXX};
assign registers[265] = {32'b01111010000000000000000011001000};
assign registers[266] = {32'b00010110001001010000100XXXXXXXXX};
assign registers[267] = {32'b01111010000000000000000000000000};
assign registers[268] = {32'b01111010100000000000000000000000};
assign registers[269] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[270] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[271] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[272] = {32'b01111011000000000000000000000010};
assign registers[273] = {32'b00010100101011011001100XXXXXXXXX};
assign registers[274] = {32'b0011XXXX0010001100XXXXXXXXXXXXXX};
assign registers[275] = {32'b10000010XXXXXXXXXX00100XXXXXXXXX};
assign registers[276] = {32'b01111010000000000000000000000000};
assign registers[277] = {32'b1000000010100XXXXX00010XXXXXXXXX};
assign registers[278] = {32'b01111010000000000000000010011101};
assign registers[279] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[280] = {32'b1000000010100XXXXX00101XXXXXXXXX};
assign registers[281] = {32'b01111010000000000000000011001000};
assign registers[282] = {32'b00010100001011010000101XXXXXXXXX};
assign registers[283] = {32'b00010100001010010000101XXXXXXXXX};
assign registers[284] = {32'b01111010000000000000000000000000};
assign registers[285] = {32'b01111010100000000000000000000000};
assign registers[286] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[287] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[288] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[289] = {32'b01000101000101010100000100100001};
assign registers[290] = {32'b01000000000000000000001000010111};
assign registers[291] = {32'b00010100001010010000110XXXXXXXXX};
assign registers[292] = {32'b01111010000000000000000000000001};
assign registers[293] = {32'b00010110001101010000110XXXXXXXXX};
assign registers[294] = {32'b01111010000000000000000000000001};
assign registers[295] = {32'b00010100000101010001101XXXXXXXXX};
assign registers[296] = {32'b01111010000000000000000000000000};
assign registers[297] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[298] = {32'b00010100101000110110100XXXXXXXXX};
assign registers[299] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[300] = {32'b010100001101110100XXXXX000000000};
assign registers[301] = {32'b00010101110111101111111111111111};
assign registers[302] = {32'b01111010000000000000000010011101};
assign registers[303] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[304] = {32'b010100001101110100XXXXX000000000};
assign registers[305] = {32'b00010101110111101111111111111111};
assign registers[306] = {32'b010100001100100010XXXXX000000000};
assign registers[307] = {32'b010100001100100011XXXXX000000001};
assign registers[308] = {32'b010100001100100100XXXXX000000010};
assign registers[309] = {32'b010100001100100101XXXXX000000011};
assign registers[310] = {32'b010100001100100110XXXXX000000100};
assign registers[311] = {32'b010100001100100111XXXXX000000101};
assign registers[312] = {32'b010100001100101000XXXXX000000110};
assign registers[313] = {32'b010100001100101001XXXXX000000111};
assign registers[314] = {32'b00010101110011100100000000001000};
assign registers[315] = {32'b010100001100101100XXXXX000000000};
assign registers[316] = {32'b010100001100101101XXXXX000000001};
assign registers[317] = {32'b00010101110011100100000000000010};
assign registers[318] = {32'b010100001100111010XXXXX000000000};
assign registers[319] = {32'b00010101110011100100000000000001};
assign registers[320] = {32'b01000001000000000000000000110011};
assign registers[321] = {32'b00010101110011100111111111111111};
assign registers[322] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[323] = {32'b00010101110011100111111111111110};
assign registers[324] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[325] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[326] = {32'b00010101110011100111111111111000};
assign registers[327] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[328] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[329] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[330] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[331] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[332] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[333] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[334] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[335] = {32'b01111010000000000000000000000000};
assign registers[336] = {32'b01111010100000000000000010011101};
assign registers[337] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[338] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[339] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[340] = {32'b010100001101110101XXXXX000000000};
assign registers[341] = {32'b00010101110111101111111111111111};
assign registers[342] = {32'b01111010000000000000000000000001};
assign registers[343] = {32'b01111010100000000000000010011101};
assign registers[344] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[345] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[346] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[347] = {32'b010100001101110101XXXXX000000000};
assign registers[348] = {32'b00010101110111101111111111111111};
assign registers[349] = {32'b010100001101100101XXXXX000000000};
assign registers[350] = {32'b00010101110111101111111111111111};
assign registers[351] = {32'b010100001100100010XXXXX000000000};
assign registers[352] = {32'b010100001100100011XXXXX000000001};
assign registers[353] = {32'b010100001100100100XXXXX000000010};
assign registers[354] = {32'b010100001100100101XXXXX000000011};
assign registers[355] = {32'b010100001100100110XXXXX000000100};
assign registers[356] = {32'b010100001100100111XXXXX000000101};
assign registers[357] = {32'b010100001100101000XXXXX000000110};
assign registers[358] = {32'b010100001100101001XXXXX000000111};
assign registers[359] = {32'b00010101110011100100000000001000};
assign registers[360] = {32'b010100001100101100XXXXX000000000};
assign registers[361] = {32'b010100001100101101XXXXX000000001};
assign registers[362] = {32'b00010101110011100100000000000010};
assign registers[363] = {32'b010100001100111010XXXXX000000000};
assign registers[364] = {32'b00010101110011100100000000000001};
assign registers[365] = {32'b01000001000000000000000000011110};
assign registers[366] = {32'b00010101110011100111111111111111};
assign registers[367] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[368] = {32'b00010101110011100111111111111110};
assign registers[369] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[370] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[371] = {32'b00010101110011100111111111111000};
assign registers[372] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[373] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[374] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[375] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[376] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[377] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[378] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[379] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[380] = {32'b1000000011000XXXXX00011XXXXXXXXX};
assign registers[381] = {32'b01111010000000000000000000000001};
assign registers[382] = {32'b00010100001011010000101XXXXXXXXX};
assign registers[383] = {32'b01111010000000000000000000000111};
assign registers[384] = {32'b0010XXXX1010000010XXXXXXXXXXXXXX};
assign registers[385] = {32'b10000010XXXXXXXXXX00111XXXXXXXXX};
assign registers[386] = {32'b01111010000000000000000000000011};
assign registers[387] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[388] = {32'b01111010100000000000000000000001};
assign registers[389] = {32'b00010100000101010110100XXXXXXXXX};
assign registers[390] = {32'b01111011000000000000000000010101};
assign registers[391] = {32'b00010100101101101010110XXXXXXXXX};
assign registers[392] = {32'b00010100101100011110111XXXXXXXXX};
assign registers[393] = {32'b010100001011110100XXXXX000000000};
assign registers[394] = {32'b01111010000000000000000000000001};
assign registers[395] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[396] = {32'b01111010000000000000000000000000};
assign registers[397] = {32'b1000000010100XXXXX10101XXXXXXXXX};
assign registers[398] = {32'b01111011000000000000000000010101};
assign registers[399] = {32'b00010100101101101010110XXXXXXXXX};
assign registers[400] = {32'b00010100101100011110111XXXXXXXXX};
assign registers[401] = {32'b010100001011110101XXXXX000000000};
assign registers[402] = {32'b01111010000000000000000000000001};
assign registers[403] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[404] = {32'b1000000000101XXXXX10100XXXXXXXXX};
assign registers[405] = {32'b01111010100000000000000000010101};
assign registers[406] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[407] = {32'b00010100101010011110110XXXXXXXXX};
assign registers[408] = {32'b010100001011010100XXXXX000000000};
assign registers[409] = {32'b01111010000000000000000000000001};
assign registers[410] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[411] = {32'b1000000000011XXXXX10100XXXXXXXXX};
assign registers[412] = {32'b01111010100000000000000000010101};
assign registers[413] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[414] = {32'b00010100101010011110110XXXXXXXXX};
assign registers[415] = {32'b010100001011010100XXXXX000000000};
assign registers[416] = {32'b01111010000000000000000000000001};
assign registers[417] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[418] = {32'b00010100001010001100101XXXXXXXXX};
assign registers[419] = {32'b1000000000101XXXXX01000XXXXXXXXX};
assign registers[420] = {32'b1000000000101XXXXX10100XXXXXXXXX};
assign registers[421] = {32'b01111010100000000000000000010101};
assign registers[422] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[423] = {32'b00010100101010011110110XXXXXXXXX};
assign registers[424] = {32'b010100001011010100XXXXX000000000};
assign registers[425] = {32'b01111010000000000000000000000001};
assign registers[426] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[427] = {32'b01111010000000000000000000101000};
assign registers[428] = {32'b00010100001011010000101XXXXXXXXX};
assign registers[429] = {32'b1000000000101XXXXX10100XXXXXXXXX};
assign registers[430] = {32'b01111010100000000000000000010101};
assign registers[431] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[432] = {32'b00010100101010011110110XXXXXXXXX};
assign registers[433] = {32'b010100001011010100XXXXX000000000};
assign registers[434] = {32'b01111010000000000000000000000001};
assign registers[435] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[436] = {32'b1000000000110XXXXX10100XXXXXXXXX};
assign registers[437] = {32'b01111010100000000000000000010101};
assign registers[438] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[439] = {32'b00010100101010011110110XXXXXXXXX};
assign registers[440] = {32'b010100001011010100XXXXX000000000};
assign registers[441] = {32'b01111010000000000000000000000111};
assign registers[442] = {32'b0010XXXX1010000010XXXXXXXXXXXXXX};
assign registers[443] = {32'b10000010XXXXXXXXXX00111XXXXXXXXX};
assign registers[444] = {32'b01111010000000000000000000000111};
assign registers[445] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[446] = {32'b01111010000000000000000000000001};
assign registers[447] = {32'b00010100001111010001000XXXXXXXXX};
assign registers[448] = {32'b01111010000000000000000000000001};
assign registers[449] = {32'b00010100010001010001001XXXXXXXXX};
assign registers[450] = {32'b01111010000000000000000000010101};
assign registers[451] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[452] = {32'b00010100101000011110100XXXXXXXXX};
assign registers[453] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[454] = {32'b010100001101110100XXXXX000000000};
assign registers[455] = {32'b00010101110111101111111111111111};
assign registers[456] = {32'b01111010000000000000000000010101};
assign registers[457] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[458] = {32'b00010100101000100010100XXXXXXXXX};
assign registers[459] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[460] = {32'b010100001101110100XXXXX000000000};
assign registers[461] = {32'b00010101110111101111111111111111};
assign registers[462] = {32'b01111010000000000000000000010101};
assign registers[463] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[464] = {32'b00010100101000100110100XXXXXXXXX};
assign registers[465] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[466] = {32'b010100001101110100XXXXX000000000};
assign registers[467] = {32'b00010101110111101111111111111111};
assign registers[468] = {32'b01111010000000000000000000000001};
assign registers[469] = {32'b00010100000101010001110XXXXXXXXX};
assign registers[470] = {32'b010100001101101110XXXXX000000000};
assign registers[471] = {32'b00010101110111101111111111111111};
assign registers[472] = {32'b010100001100100010XXXXX000000000};
assign registers[473] = {32'b010100001100100011XXXXX000000001};
assign registers[474] = {32'b010100001100100100XXXXX000000010};
assign registers[475] = {32'b010100001100100101XXXXX000000011};
assign registers[476] = {32'b010100001100100110XXXXX000000100};
assign registers[477] = {32'b010100001100100111XXXXX000000101};
assign registers[478] = {32'b010100001100101000XXXXX000000110};
assign registers[479] = {32'b010100001100101001XXXXX000000111};
assign registers[480] = {32'b00010101110011100100000000001000};
assign registers[481] = {32'b010100001100101100XXXXX000000000};
assign registers[482] = {32'b010100001100101101XXXXX000000001};
assign registers[483] = {32'b010100001100101110XXXXX000000010};
assign registers[484] = {32'b00010101110011100100000000000011};
assign registers[485] = {32'b010100001100111010XXXXX000000000};
assign registers[486] = {32'b00010101110011100100000000000001};
assign registers[487] = {32'b01000001000000000000000000111111};
assign registers[488] = {32'b00010101110011100111111111111111};
assign registers[489] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[490] = {32'b00010101110011100111111111111101};
assign registers[491] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[492] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[493] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[494] = {32'b00010101110011100111111111111000};
assign registers[495] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[496] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[497] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[498] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[499] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[500] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[501] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[502] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[503] = {32'b01111010000000000000000000000001};
assign registers[504] = {32'b00010100000101010000010XXXXXXXXX};
assign registers[505] = {32'b01111010000000000000000000000001};
assign registers[506] = {32'b00010100001101010000110XXXXXXXXX};
assign registers[507] = {32'b1000000000110XXXXX00101XXXXXXXXX};
assign registers[508] = {32'b01111010000000000000000000000001};
assign registers[509] = {32'b01111010100000000000000000010101};
assign registers[510] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[511] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[512] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[513] = {32'b1000000010101XXXXX00111XXXXXXXXX};
assign registers[514] = {32'b01111010000000000000000000000001};
assign registers[515] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[516] = {32'b1000000000111XXXXX10100XXXXXXXXX};
assign registers[517] = {32'b01111010100000000000000000010101};
assign registers[518] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[519] = {32'b01111011000000000000000000000001};
assign registers[520] = {32'b00010100101011011010110XXXXXXXXX};
assign registers[521] = {32'b010100001011010100XXXXX000000000};
assign registers[522] = {32'b01111010000000000000000000000010};
assign registers[523] = {32'b01111010100000000000000000010101};
assign registers[524] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[525] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[526] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[527] = {32'b1000000010101XXXXX00111XXXXXXXXX};
assign registers[528] = {32'b01111010000000000000000000000001};
assign registers[529] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[530] = {32'b1000000000111XXXXX10100XXXXXXXXX};
assign registers[531] = {32'b01111010100000000000000000010101};
assign registers[532] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[533] = {32'b01111011000000000000000000000010};
assign registers[534] = {32'b00010100101011011010110XXXXXXXXX};
assign registers[535] = {32'b010100001011010100XXXXX000000000};
assign registers[536] = {32'b01000000000000000000000100011010};
assign registers[537] = {32'b01111010000000000000000000000000};
assign registers[538] = {32'b01111010100000000000000000010101};
assign registers[539] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[540] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[541] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[542] = {32'b1000000010101XXXXX00111XXXXXXXXX};
assign registers[543] = {32'b01111010000000000000000000000001};
assign registers[544] = {32'b00010110001111010000111XXXXXXXXX};
assign registers[545] = {32'b1000000000111XXXXX10100XXXXXXXXX};
assign registers[546] = {32'b01111010100000000000000000010101};
assign registers[547] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[548] = {32'b01111011000000000000000000000000};
assign registers[549] = {32'b00010100101011011010110XXXXXXXXX};
assign registers[550] = {32'b010100001011010100XXXXX000000000};
assign registers[551] = {32'b01111010000000000000000000000000};
assign registers[552] = {32'b01111010100000000000000000010101};
assign registers[553] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[554] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[555] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[556] = {32'b1000000010101XXXXX00010XXXXXXXXX};
assign registers[557] = {32'b01111010000000000000000000000001};
assign registers[558] = {32'b00010100000101010000010XXXXXXXXX};
assign registers[559] = {32'b01111010000000000000000000000010};
assign registers[560] = {32'b01111010100000000000000000010101};
assign registers[561] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[562] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[563] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[564] = {32'b01001000000101010100001000110100};
assign registers[565] = {32'b01000000000000000000001000110110};
assign registers[566] = {32'b01111010000000000000000000000000};
assign registers[567] = {32'b1000000010100XXXXX00010XXXXXXXXX};
assign registers[568] = {32'b01111010000000000000000000000111};
assign registers[569] = {32'b0010XXXX1010000010XXXXXXXXXXXXXX};
assign registers[570] = {32'b10000010XXXXXXXXXX00111XXXXXXXXX};
assign registers[571] = {32'b01111010000000000000000000000100};
assign registers[572] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[573] = {32'b01111010000000000000000000010101};
assign registers[574] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[575] = {32'b00010100101000011110100XXXXXXXXX};
assign registers[576] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[577] = {32'b01111010100000000000000000000000};
assign registers[578] = {32'b01000100101001010100001001000010};
assign registers[579] = {32'b01000000000000000000001001010010};
assign registers[580] = {32'b01111010000000000000000000000001};
assign registers[581] = {32'b00010100000101010000010XXXXXXXXX};
assign registers[582] = {32'b01111010000000000000000000000111};
assign registers[583] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[584] = {32'b01111010000000000000000000000010};
assign registers[585] = {32'b01111010100000000000000000010101};
assign registers[586] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[587] = {32'b00010100101011010010101XXXXXXXXX};
assign registers[588] = {32'b0110XXXX10101XXXXX10101000000000};
assign registers[589] = {32'b01001000000101010100001001001101};
assign registers[590] = {32'b01000000000000000000001001010001};
assign registers[591] = {32'b01111010000000000000000000000000};
assign registers[592] = {32'b1000000010100XXXXX00010XXXXXXXXX};
assign registers[593] = {32'b01111010000000000000000000000100};
assign registers[594] = {32'b1000000010100XXXXX00111XXXXXXXXX};
assign registers[595] = {32'b01000000000000000000001000111011};
assign registers[596] = {32'b010100001101100010XXXXX000000000};
assign registers[597] = {32'b00010101110111101111111111111111};
assign registers[598] = {32'b010100001100100010XXXXX000000000};
assign registers[599] = {32'b010100001100100011XXXXX000000001};
assign registers[600] = {32'b010100001100100100XXXXX000000010};
assign registers[601] = {32'b010100001100100101XXXXX000000011};
assign registers[602] = {32'b010100001100100110XXXXX000000100};
assign registers[603] = {32'b010100001100100111XXXXX000000101};
assign registers[604] = {32'b010100001100101000XXXXX000000110};
assign registers[605] = {32'b010100001100101001XXXXX000000111};
assign registers[606] = {32'b00010101110011100100000000001000};
assign registers[607] = {32'b010100001100101100XXXXX000000000};
assign registers[608] = {32'b010100001100101101XXXXX000000001};
assign registers[609] = {32'b010100001100101110XXXXX000000010};
assign registers[610] = {32'b00010101110011100100000000000011};
assign registers[611] = {32'b010100001100111010XXXXX000000000};
assign registers[612] = {32'b00010101110011100100000000000001};
assign registers[613] = {32'b01000001000000000000000000010100};
assign registers[614] = {32'b00010101110011100111111111111111};
assign registers[615] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[616] = {32'b00010101110011100111111111111101};
assign registers[617] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[618] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[619] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[620] = {32'b00010101110011100111111111111000};
assign registers[621] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[622] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[623] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[624] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[625] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[626] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[627] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[628] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[629] = {32'b1000000000010XXXXX10100XXXXXXXXX};
assign registers[630] = {32'b01111010100000000000000000010101};
assign registers[631] = {32'b00010100101011101010101XXXXXXXXX};
assign registers[632] = {32'b01111011000000000000000000000000};
assign registers[633] = {32'b00010100101011011010110XXXXXXXXX};
assign registers[634] = {32'b010100001011010100XXXXX000000000};
assign registers[635] = {32'b01111010000000000000000000000111};
assign registers[636] = {32'b0010XXXX1010000010XXXXXXXXXXXXXX};
assign registers[637] = {32'b10000010XXXXXXXXXX00111XXXXXXXXX};
assign registers[638] = {32'b01111010000000000000000000000101};
assign registers[639] = {32'b00010100001111010000111XXXXXXXXX};
assign registers[640] = {32'b01111010000000000000000000000001};
assign registers[641] = {32'b00010100001111010001000XXXXXXXXX};
assign registers[642] = {32'b01111010000000000000000000000001};
assign registers[643] = {32'b00010100010001010001001XXXXXXXXX};
assign registers[644] = {32'b01111010000000000000000000010101};
assign registers[645] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[646] = {32'b00010100101000011110100XXXXXXXXX};
assign registers[647] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[648] = {32'b010100001101110100XXXXX000000000};
assign registers[649] = {32'b00010101110111101111111111111111};
assign registers[650] = {32'b01111010000000000000000000010101};
assign registers[651] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[652] = {32'b00010100101000100010100XXXXXXXXX};
assign registers[653] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[654] = {32'b010100001101110100XXXXX000000000};
assign registers[655] = {32'b00010101110111101111111111111111};
assign registers[656] = {32'b01111010000000000000000000010101};
assign registers[657] = {32'b00010100101001101010100XXXXXXXXX};
assign registers[658] = {32'b00010100101000100110100XXXXXXXXX};
assign registers[659] = {32'b0110XXXX10100XXXXX10100000000000};
assign registers[660] = {32'b010100001101110100XXXXX000000000};
assign registers[661] = {32'b00010101110111101111111111111111};
assign registers[662] = {32'b010100001100100010XXXXX000000000};
assign registers[663] = {32'b010100001100100011XXXXX000000001};
assign registers[664] = {32'b010100001100100100XXXXX000000010};
assign registers[665] = {32'b010100001100100101XXXXX000000011};
assign registers[666] = {32'b010100001100100110XXXXX000000100};
assign registers[667] = {32'b010100001100100111XXXXX000000101};
assign registers[668] = {32'b010100001100101000XXXXX000000110};
assign registers[669] = {32'b010100001100101001XXXXX000000111};
assign registers[670] = {32'b00010101110011100100000000001000};
assign registers[671] = {32'b010100001100101100XXXXX000000000};
assign registers[672] = {32'b010100001100101101XXXXX000000001};
assign registers[673] = {32'b010100001100101110XXXXX000000010};
assign registers[674] = {32'b00010101110011100100000000000011};
assign registers[675] = {32'b010100001100111010XXXXX000000000};
assign registers[676] = {32'b00010101110011100100000000000001};
assign registers[677] = {32'b01000001000000000000000001100100};
assign registers[678] = {32'b00010101110011100111111111111111};
assign registers[679] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[680] = {32'b00010101110011100111111111111101};
assign registers[681] = {32'b0110XXXX11001XXXXX01100000000000};
assign registers[682] = {32'b0110XXXX11001XXXXX01101000000001};
assign registers[683] = {32'b0110XXXX11001XXXXX01110000000010};
assign registers[684] = {32'b00010101110011100111111111111000};
assign registers[685] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[686] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[687] = {32'b0110XXXX11001XXXXX00100000000010};
assign registers[688] = {32'b0110XXXX11001XXXXX00101000000011};
assign registers[689] = {32'b0110XXXX11001XXXXX00110000000100};
assign registers[690] = {32'b0110XXXX11001XXXXX00111000000101};
assign registers[691] = {32'b0110XXXX11001XXXXX01000000000110};
assign registers[692] = {32'b0110XXXX11001XXXXX01001000000111};
assign registers[693] = {32'b10110010XXXXXXXXXXXXXXXXXXXXXXXX};
assign registers[694] = {32'b00000001000000000000000000000000};
assign registers[695] = {32'b11111111111111111111111111111111};

//Meus arquivos de programas que serao executados
assign registers[4096] = {16'd0, 16'd4};
//Programa 1 estara na track 2 no setor 0
assign registers[4097] = {16'd0, 8'd2, 8'd0};
//Programa 2 estara na track 2 no setor 1
assign registers[4098] = {16'd0, 8'd2, 8'd1};
assign registers[4099] = {32'b11111111111111111111111111111111};
//Fim dos arquivos de programas

//Programa teste 1 
assign registers[8192] = {16'd0, 16'd33};
assign registers[8193] = {32'b01110000000000000000000000000000};
assign registers[8194] = {32'b01000000000000000000000000001001};
assign registers[8195] = {32'b0110XXXX11010XXXXX11001111111110};
assign registers[8196] = {32'b0110XXXX11010XXXXX10100111111111};
assign registers[8197] = {32'b0100001010100XXXXXXXXXXXXXXXXXXX};
assign registers[8198] = {32'b00010101110111101100000000000001};
assign registers[8199] = {32'b0110XXXX11011XXXXX01101000000000};
assign registers[8200] = {32'b1010XXXX0110100000XXXX0000000000};
assign registers[8201] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[8202] = {32'b1000000011001XXXXX11010XXXXXXXXX};
assign registers[8203] = {32'b01111010000000000000000000000010};
assign registers[8204] = {32'b1000000010100XXXXX00010XXXXXXXXX};
assign registers[8205] = {32'b01111010000000000000000000000001};
assign registers[8206] = {32'b01111010100000000000000000000001};
assign registers[8207] = {32'b01000011101001010100000000010000};
assign registers[8208] = {32'b01000000000000000000000000011110};
assign registers[8209] = {32'b010100001101100010XXXXX000000000};
assign registers[8210] = {32'b00010101110111101111111111111111};
assign registers[8211] = {32'b010100001100100010XXXXX000000000};
assign registers[8212] = {32'b00010101110011100100000000000001};
assign registers[8213] = {32'b010100001100111010XXXXX000000000};
assign registers[8214] = {32'b00010101110011100100000000000001};
assign registers[8215] = {32'b01000001000000000000000000000101};
assign registers[8216] = {32'b00010101110011100111111111111111};
assign registers[8217] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[8218] = {32'b00010101110011100111111111111111};
assign registers[8219] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[8220] = {32'b01111010000000000000000000000010};
assign registers[8221] = {32'b00010100000101010000010XXXXXXXXX};
assign registers[8222] = {32'b01000000000000000000000000001100};
assign registers[8223] = {32'b00000001000000000000000000000000};
assign registers[8224] = {32'b11111111111111111111111111111111};

//Programa teste 2
assign registers[8320] = {16'd0, 16'd38};
assign registers[8321] = {32'b01110000000000000000000000000000};
assign registers[8322] = {32'b01000000000000000000000000001001};
assign registers[8323] = {32'b0110XXXX11010XXXXX11001111111110};
assign registers[8324] = {32'b0110XXXX11010XXXXX10100111111111};
assign registers[8325] = {32'b0100001010100XXXXXXXXXXXXXXXXXXX};
assign registers[8326] = {32'b00010101110111101100000000000001};
assign registers[8327] = {32'b0110XXXX11011XXXXX01101000000000};
assign registers[8328] = {32'b1010XXXX0110100000XXXX0000000000};
assign registers[8329] = {32'b0100001011111XXXXXXXXXXXXXXXXXXX};
assign registers[8330] = {32'b1000000011001XXXXX11010XXXXXXXXX};
assign registers[8331] = {32'b01111010000000000000000000000000};
assign registers[8332] = {32'b1000000010100XXXXX00010XXXXXXXXX};
assign registers[8333] = {32'b01111010000000000000000000001011};
assign registers[8334] = {32'b1000000010100XXXXX00011XXXXXXXXX};
assign registers[8335] = {32'b01111010000000000000000000000010};
assign registers[8336] = {32'b01000101000101010000000000010001};
assign registers[8337] = {32'b01000000000000000000000000100011};
assign registers[8338] = {32'b010100001101100011XXXXX000000000};
assign registers[8339] = {32'b00010101110111101111111111111111};
assign registers[8340] = {32'b010100001100100010XXXXX000000000};
assign registers[8341] = {32'b010100001100100011XXXXX000000001};
assign registers[8342] = {32'b00010101110011100100000000000010};
assign registers[8343] = {32'b010100001100111010XXXXX000000000};
assign registers[8344] = {32'b00010101110011100100000000000001};
assign registers[8345] = {32'b01000001000000000000000000000101};
assign registers[8346] = {32'b00010101110011100111111111111111};
assign registers[8347] = {32'b0110XXXX11001XXXXX11010000000000};
assign registers[8348] = {32'b00010101110011100111111111111110};
assign registers[8349] = {32'b0110XXXX11001XXXXX00010000000000};
assign registers[8350] = {32'b0110XXXX11001XXXXX00011000000001};
assign registers[8351] = {32'b01111010000000000000000000000001};
assign registers[8352] = {32'b00010100000101010000010XXXXXXXXX};
assign registers[8353] = {32'b01111010000000000000000000000010};
assign registers[8354] = {32'b00010100000111010000011XXXXXXXXX};
assign registers[8355] = {32'b01000000000000000000000000001110};
assign registers[8356] = {32'b00000001000000000000000000000000};
assign registers[8357] = {32'b11111111111111111111111111111111};

endmodule 